VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tiny_user_project
  CLASS BLOCK ;
  FOREIGN tiny_user_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 981.120 1.000 981.680 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 1.000 57.680 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 450.240 999.000 450.800 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 215.040 4.000 215.600 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 996.000 323.120 999.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 658.560 999.000 659.120 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 996.000 272.720 999.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 104.160 4.000 104.720 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 957.600 999.000 958.160 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 336.000 4.000 336.560 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 996.000 356.720 999.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 1.000 91.280 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 996.000 239.120 999.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 996.000 289.520 999.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 90.720 4.000 91.280 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 248.640 4.000 249.200 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 745.920 999.000 746.480 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 996.000 20.720 999.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 996.000 622.160 999.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 996.000 259.280 999.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 36.960 4.000 37.520 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 996.000 444.080 999.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 816.480 4.000 817.040 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 1.000 427.280 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 288.960 4.000 289.520 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 996.000 672.560 999.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 996.000 575.120 999.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 1.000 302.960 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 665.280 999.000 665.840 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 342.720 4.000 343.280 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 927.360 1.000 927.920 4.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 349.440 4.000 350.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 944.160 996.000 944.720 999.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 131.040 999.000 131.600 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 594.720 999.000 595.280 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 551.040 4.000 551.600 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 467.040 996.000 467.600 999.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 645.120 4.000 645.680 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 362.880 999.000 363.440 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 342.720 999.000 343.280 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 996.000 588.560 999.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 996.000 336.560 999.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 742.560 1.000 743.120 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 996.000 158.480 999.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 369.600 999.000 370.160 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 685.440 1.000 686.000 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 987.840 4.000 988.400 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 996.000 7.280 999.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 302.400 4.000 302.960 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 1.000 679.280 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 996.000 165.200 999.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 996.000 679.280 999.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 178.080 4.000 178.640 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 416.640 999.000 417.200 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 991.200 999.000 991.760 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 776.160 4.000 776.720 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 996.000 98.000 999.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 10.080 4.000 10.640 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 601.440 996.000 602.000 999.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 739.200 999.000 739.760 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 863.520 999.000 864.080 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 1.000 625.520 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 876.960 4.000 877.520 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 996.000 111.440 999.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 996.000 27.440 999.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 996.000 171.920 999.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 540.960 4.000 541.520 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 1.000 447.440 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 729.120 4.000 729.680 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 996.000 759.920 999.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 1.000 507.920 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 268.800 4.000 269.360 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 712.320 996.000 712.880 999.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 964.320 996.000 964.880 999.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 705.600 4.000 706.160 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 996.000 87.920 999.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 974.400 4.000 974.960 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 937.440 996.000 938.000 999.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 453.600 4.000 454.160 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 930.720 999.000 931.280 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 322.560 4.000 323.120 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 1.000 131.600 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 779.520 999.000 780.080 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 238.560 999.000 239.120 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 651.840 999.000 652.400 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 897.120 999.000 897.680 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 786.240 999.000 786.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 1.000 118.160 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 769.440 1.000 770.000 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 960.960 4.000 961.520 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 954.240 1.000 954.800 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 1.000 558.320 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 117.600 999.000 118.160 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 678.720 4.000 679.280 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 996.000 185.360 999.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 6.720 999.000 7.280 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 561.120 999.000 561.680 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 1.000 235.760 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 957.600 996.000 958.160 999.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 1.000 316.400 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 883.680 999.000 884.240 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 907.200 1.000 907.760 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 759.360 999.000 759.920 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 991.200 996.000 991.760 999.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 678.720 999.000 679.280 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 996.000 178.640 999.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 903.840 1.000 904.400 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 487.200 4.000 487.760 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 104.160 999.000 104.720 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 628.320 999.000 628.880 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 996.000 494.480 999.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 228.480 4.000 229.040 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 996.000 397.040 999.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 967.680 4.000 968.240 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 1.000 323.120 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 409.920 999.000 410.480 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 786.240 996.000 786.800 999.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 514.080 999.000 514.640 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 288.960 999.000 289.520 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.080 996.000 430.640 999.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 996.000 145.040 999.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 917.280 999.000 917.840 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 749.280 4.000 749.840 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 635.040 999.000 635.600 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 110.880 999.000 111.440 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 996.000 534.800 999.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 272.160 999.000 272.720 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 996.000 706.160 999.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 769.440 4.000 770.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 1.000 30.800 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 638.400 999.000 638.960 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 782.880 4.000 783.440 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 164.640 999.000 165.200 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 732.480 996.000 733.040 999.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 1.000 242.480 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 1.000 440.720 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 996.000 390.320 999.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 799.680 996.000 800.240 999.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 608.160 999.000 608.720 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 719.040 4.000 719.600 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 996.000 665.840 999.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 974.400 1.000 974.960 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 996.000 34.160 999.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 20.160 999.000 20.720 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 996.000 74.480 999.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 255.360 4.000 255.920 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 762.720 1.000 763.280 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 534.240 4.000 534.800 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 446.880 4.000 447.440 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 890.400 1.000 890.960 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 725.760 999.000 726.320 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 157.920 4.000 158.480 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 430.080 999.000 430.640 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 406.560 4.000 407.120 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 843.360 999.000 843.920 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 752.640 996.000 753.200 999.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 1.000 249.200 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 996.000 0.560 999.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 30.240 4.000 30.800 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 1.000 665.840 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 534.240 999.000 534.800 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 204.960 999.000 205.520 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 658.560 4.000 659.120 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 806.400 999.000 806.960 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 70.560 4.000 71.120 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 601.440 999.000 602.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 1.000 719.600 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 796.320 1.000 796.880 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 940.800 1.000 941.360 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 996.000 350.000 999.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 729.120 1.000 729.680 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 1.000 413.840 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 996.000 450.800 999.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 829.920 4.000 830.480 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 779.520 996.000 780.080 999.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 971.040 996.000 971.600 999.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 443.520 999.000 444.080 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 1.000 17.360 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 514.080 4.000 514.640 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 1.000 202.160 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 1.000 262.640 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 460.320 999.000 460.880 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 772.800 999.000 773.360 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 996.000 316.400 999.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 171.360 4.000 171.920 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 544.320 4.000 544.880 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 1.000 672.560 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 698.880 996.000 699.440 999.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 1.000 195.440 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 1.000 350.000 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 16.800 4.000 17.360 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 994.560 4.000 995.120 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 950.880 996.000 951.440 999.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 198.240 999.000 198.800 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 1.000 124.880 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 1.000 474.320 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 1.000 3.920 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 749.280 1.000 749.840 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 823.200 996.000 823.760 999.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 876.960 1.000 877.520 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 420.000 4.000 420.560 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 996.000 61.040 999.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 1.000 208.880 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 252.000 999.000 252.560 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 557.760 4.000 558.320 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 944.160 999.000 944.720 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 1.000 870.800 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 934.080 4.000 934.640 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 996.000 403.760 999.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 241.920 4.000 242.480 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 732.480 999.000 733.040 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 403.200 999.000 403.760 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 258.720 999.000 259.280 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 191.520 999.000 192.080 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 996.000 232.400 999.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 994.560 1.000 995.120 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 1.000 494.480 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 1.000 393.680 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 1.000 487.760 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 645.120 999.000 645.680 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 799.680 999.000 800.240 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 282.240 999.000 282.800 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 315.840 999.000 316.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 823.200 1.000 823.760 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 322.560 999.000 323.120 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 440.160 4.000 440.720 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 996.000 830.480 999.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 3.360 4.000 3.920 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 996.000 383.600 999.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 712.320 999.000 712.880 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 500.640 4.000 501.200 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 604.800 4.000 605.360 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 996.000 329.840 999.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 996.000 218.960 999.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 996.000 568.400 999.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 996.000 14.000 999.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 26.880 999.000 27.440 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 1.000 356.720 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 1.000 400.400 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 90.720 999.000 91.280 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 356.160 4.000 356.720 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 870.240 4.000 870.800 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 473.760 999.000 474.320 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 672.000 4.000 672.560 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 1.000 178.640 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 624.960 4.000 625.520 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 924.000 996.000 924.560 999.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 863.520 4.000 864.080 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 84.000 4.000 84.560 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 376.320 999.000 376.880 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 547.680 999.000 548.240 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 315.840 4.000 316.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 996.000 212.240 999.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 658.560 1.000 659.120 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 789.600 4.000 790.160 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 996.000 507.920 999.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 996.000 595.280 999.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 1.000 158.480 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 725.760 996.000 726.320 999.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 903.840 996.000 904.400 999.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 77.280 4.000 77.840 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 996.000 410.480 999.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 876.960 999.000 877.520 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 231.840 999.000 232.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 235.200 4.000 235.760 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 1.000 380.240 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 362.880 4.000 363.440 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 1.000 571.760 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 40.320 999.000 40.880 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 996.000 151.760 999.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 917.280 996.000 917.840 999.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 796.320 4.000 796.880 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 329.280 4.000 329.840 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 913.920 1.000 914.480 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 577.920 1.000 578.480 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 598.080 4.000 598.640 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 890.400 999.000 890.960 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 453.600 999.000 454.160 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 386.400 4.000 386.960 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 500.640 999.000 501.200 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 987.840 1.000 988.400 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 996.000 67.760 999.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 178.080 999.000 178.640 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 638.400 4.000 638.960 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 996.000 54.320 999.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 971.040 999.000 971.600 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 201.600 4.000 202.160 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 645.120 996.000 645.680 999.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 383.040 999.000 383.600 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 1.000 460.880 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 996.000 548.240 999.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 194.880 4.000 195.440 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 467.040 999.000 467.600 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 1.000 151.760 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 920.640 4.000 921.200 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 151.200 999.000 151.760 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 467.040 1.000 467.600 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 295.680 4.000 296.240 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 996.000 198.800 999.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 996.000 561.680 999.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 967.680 1.000 968.240 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 876.960 996.000 877.520 999.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 742.560 4.000 743.120 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 473.760 4.000 474.320 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 792.960 996.000 793.520 999.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 275.520 999.000 276.080 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 996.000 370.160 999.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 631.680 4.000 632.240 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 564.480 1.000 565.040 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 996.000 296.240 999.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 996.000 266.000 999.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 843.360 1.000 843.920 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 33.600 999.000 34.160 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 984.480 996.000 985.040 999.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 996.000 343.280 999.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 117.600 4.000 118.160 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 1.000 71.120 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 467.040 4.000 467.600 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 564.480 4.000 565.040 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 1.000 309.680 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 756.000 4.000 756.560 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 507.360 999.000 507.920 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 611.520 4.000 612.080 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 480.480 999.000 481.040 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 50.400 4.000 50.960 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 1.000 528.080 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 930.720 996.000 931.280 999.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 766.080 996.000 766.640 999.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 996.000 474.320 999.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 1.000 138.320 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 1.000 790.160 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 850.080 4.000 850.640 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 540.960 999.000 541.520 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 225.120 999.000 225.680 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 137.760 999.000 138.320 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 1.000 481.040 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 712.320 1.000 712.880 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 1.000 366.800 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 897.120 996.000 897.680 999.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 1.000 544.880 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 996.000 376.880 999.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 940.800 4.000 941.360 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 1.000 269.360 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 996.000 487.760 999.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 1.000 501.200 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 97.440 999.000 98.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 947.520 1.000 948.080 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 218.400 999.000 218.960 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 171.360 999.000 171.920 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 1.000 373.520 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 913.920 4.000 914.480 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 124.320 4.000 124.880 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 996.000 205.520 999.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 816.480 1.000 817.040 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 996.000 131.600 999.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 181.440 4.000 182.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 0.000 999.000 0.560 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 520.800 999.000 521.360 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 540.960 996.000 541.520 999.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 1.000 638.960 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 996.000 514.640 999.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 996.000 521.360 999.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 756.000 1.000 756.560 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 850.080 1.000 850.640 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 843.360 996.000 843.920 999.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 996.000 309.680 999.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 996.000 417.200 999.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 782.880 1.000 783.440 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 996.000 81.200 999.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 372.960 4.000 373.520 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 816.480 996.000 817.040 999.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 13.440 999.000 14.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 1.000 454.160 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 1.000 534.800 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 984.480 999.000 985.040 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 836.640 4.000 837.200 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 836.640 996.000 837.200 999.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 1.000 255.920 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 581.280 999.000 581.840 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 996.000 454.160 999.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 977.760 996.000 978.320 999.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 567.840 999.000 568.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 651.840 996.000 652.400 999.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 772.800 996.000 773.360 999.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 1.000 407.120 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 766.080 999.000 766.640 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 735.840 1.000 736.400 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 520.800 4.000 521.360 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 1.000 188.720 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 996.000 581.840 999.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 1.000 585.200 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 1.000 521.360 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 950.880 999.000 951.440 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 396.480 999.000 397.040 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 480.480 4.000 481.040 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 574.560 999.000 575.120 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 645.120 1.000 645.680 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 1.000 363.440 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 725.760 4.000 726.320 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 829.920 999.000 830.480 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 577.920 4.000 578.480 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 685.440 4.000 686.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 1.000 830.480 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 265.440 999.000 266.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 692.160 999.000 692.720 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 164.640 4.000 165.200 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 137.760 4.000 138.320 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 540.960 1.000 541.520 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 1.000 289.520 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 184.800 999.000 185.360 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 1.000 64.400 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 1.000 296.240 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 157.920 999.000 158.480 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 937.440 999.000 938.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 423.360 999.000 423.920 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 1.000 104.720 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 309.120 4.000 309.680 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 1.000 706.160 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 996.000 870.800 999.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 651.840 1.000 652.400 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 554.400 999.000 554.960 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 997.920 996.000 998.480 999.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 883.680 996.000 884.240 999.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 43.680 4.000 44.240 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 460.320 4.000 460.880 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 996.000 276.080 999.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 1.000 336.560 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 996.000 104.720 999.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 329.280 999.000 329.840 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 588.000 999.000 588.560 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 131.040 4.000 131.600 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 1.000 776.720 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 816.480 999.000 817.040 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 665.280 4.000 665.840 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 910.560 996.000 911.120 999.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 856.800 4.000 857.360 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 934.080 1.000 934.640 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 996.000 40.880 999.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 843.360 4.000 843.920 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 73.920 999.000 74.480 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 1.000 182.000 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 1.000 276.080 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 960.960 1.000 961.520 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 309.120 999.000 309.680 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 823.200 999.000 823.760 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 692.160 4.000 692.720 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 996.000 460.880 999.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 996.000 302.960 999.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 493.920 4.000 494.480 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 924.000 999.000 924.560 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 735.840 4.000 736.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 996.000 245.840 999.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 144.480 4.000 145.040 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 813.120 999.000 813.680 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 996.000 692.720 999.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 927.360 4.000 927.920 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 806.400 996.000 806.960 999.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 856.800 996.000 857.360 999.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 863.520 996.000 864.080 999.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 1.000 598.640 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 996.000 528.080 999.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 1.000 37.520 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 1.000 10.640 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 897.120 1.000 897.680 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 413.280 4.000 413.840 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 211.680 999.000 212.240 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 527.520 4.000 528.080 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 698.880 4.000 699.440 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 954.240 4.000 954.800 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 433.440 4.000 434.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 366.240 4.000 366.800 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 282.240 4.000 282.800 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 996.000 501.200 999.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 920.640 1.000 921.200 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 1.000 434.000 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 809.760 4.000 810.320 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 698.880 999.000 699.440 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 910.560 999.000 911.120 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 584.640 4.000 585.200 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 712.320 4.000 712.880 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 124.320 999.000 124.880 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 856.800 999.000 857.360 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 996.000 363.440 999.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 719.040 999.000 719.600 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 863.520 1.000 864.080 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 507.360 4.000 507.920 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 245.280 999.000 245.840 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 996.000 282.800 999.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 47.040 999.000 47.600 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 903.840 4.000 904.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 1.000 145.040 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 379.680 4.000 380.240 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 631.680 1.000 632.240 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 850.080 999.000 850.640 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 1.000 282.800 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 60.480 999.000 61.040 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 981.120 4.000 981.680 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 614.880 996.000 615.440 999.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 151.200 4.000 151.760 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 947.520 4.000 948.080 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 996.000 47.600 999.000 ;
    END
  END la_oenb[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 984.220 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 984.220 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 302.400 999.000 302.960 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 890.400 4.000 890.960 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 275.520 4.000 276.080 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 996.000 423.920 999.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 996.000 192.080 999.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 762.720 4.000 763.280 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 1.000 98.000 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 591.360 4.000 591.920 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 903.840 999.000 904.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 836.640 999.000 837.200 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 698.880 1.000 699.440 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 63.840 4.000 64.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 436.800 999.000 437.360 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 53.760 999.000 54.320 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 996.000 437.360 999.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 745.920 996.000 746.480 999.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.240 1.000 618.800 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 883.680 1.000 884.240 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 336.000 999.000 336.560 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 883.680 4.000 884.240 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 591.360 1.000 591.920 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 1.000 111.440 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 996.000 124.880 999.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 705.600 999.000 706.160 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 890.400 996.000 890.960 999.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 1.000 420.560 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 628.320 996.000 628.880 999.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 527.520 999.000 528.080 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 836.640 1.000 837.200 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 996.000 608.720 999.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 803.040 1.000 803.600 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 1.000 343.280 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 1.000 50.960 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 67.200 999.000 67.760 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 356.160 999.000 356.720 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 996.000 138.320 999.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 997.920 999.000 998.480 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 571.200 4.000 571.760 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 651.840 4.000 652.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 97.440 4.000 98.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 1.000 44.240 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 1.000 229.040 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 614.880 999.000 615.440 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 604.800 1.000 605.360 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 996.000 554.960 999.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 813.120 996.000 813.680 999.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 897.120 4.000 897.680 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 1.000 165.200 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 685.440 999.000 686.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 850.080 996.000 850.640 999.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 426.720 4.000 427.280 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 870.240 999.000 870.800 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 389.760 999.000 390.320 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 23.520 4.000 24.080 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 739.200 996.000 739.760 999.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 996.000 118.160 999.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 1.000 329.840 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 672.000 999.000 672.560 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 856.800 1.000 857.360 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 349.440 999.000 350.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 393.120 4.000 393.680 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 80.640 999.000 81.200 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 1.000 171.920 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 1.000 514.640 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 487.200 999.000 487.760 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 996.000 719.600 999.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 964.320 999.000 964.880 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 87.360 999.000 87.920 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 1.000 84.560 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 621.600 999.000 622.160 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 1.000 24.080 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 977.760 999.000 978.320 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 685.440 996.000 686.000 999.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 144.480 999.000 145.040 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 110.880 4.000 111.440 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 188.160 4.000 188.720 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 221.760 4.000 222.320 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 1.000 692.720 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 809.760 1.000 810.320 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 399.840 4.000 400.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 803.040 4.000 803.600 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 996.000 225.680 999.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 262.080 4.000 262.640 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 1.000 215.600 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 1.000 77.840 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 996.000 481.040 999.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 996.000 252.560 999.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 1.000 551.600 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 658.560 996.000 659.120 999.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 295.680 999.000 296.240 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 618.240 4.000 618.800 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 792.960 999.000 793.520 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 1.000 222.320 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 1.000 386.960 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 57.120 4.000 57.680 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 752.640 999.000 753.200 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 1.000 612.080 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 996.000 638.960 999.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 635.040 996.000 635.600 999.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 907.200 4.000 907.760 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 996.000 91.280 999.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 725.760 1.000 726.320 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 208.320 4.000 208.880 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 823.200 4.000 823.760 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 493.920 999.000 494.480 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 992.880 984.220 ;
      LAYER Metal2 ;
        RECT 0.860 995.700 6.420 996.000 ;
        RECT 7.580 995.700 13.140 996.000 ;
        RECT 14.300 995.700 19.860 996.000 ;
        RECT 21.020 995.700 26.580 996.000 ;
        RECT 27.740 995.700 33.300 996.000 ;
        RECT 34.460 995.700 40.020 996.000 ;
        RECT 41.180 995.700 46.740 996.000 ;
        RECT 47.900 995.700 53.460 996.000 ;
        RECT 54.620 995.700 60.180 996.000 ;
        RECT 61.340 995.700 66.900 996.000 ;
        RECT 68.060 995.700 73.620 996.000 ;
        RECT 74.780 995.700 80.340 996.000 ;
        RECT 81.500 995.700 87.060 996.000 ;
        RECT 88.220 995.700 90.420 996.000 ;
        RECT 91.580 995.700 97.140 996.000 ;
        RECT 98.300 995.700 103.860 996.000 ;
        RECT 105.020 995.700 110.580 996.000 ;
        RECT 111.740 995.700 117.300 996.000 ;
        RECT 118.460 995.700 124.020 996.000 ;
        RECT 125.180 995.700 130.740 996.000 ;
        RECT 131.900 995.700 137.460 996.000 ;
        RECT 138.620 995.700 144.180 996.000 ;
        RECT 145.340 995.700 150.900 996.000 ;
        RECT 152.060 995.700 157.620 996.000 ;
        RECT 158.780 995.700 164.340 996.000 ;
        RECT 165.500 995.700 171.060 996.000 ;
        RECT 172.220 995.700 177.780 996.000 ;
        RECT 178.940 995.700 184.500 996.000 ;
        RECT 185.660 995.700 191.220 996.000 ;
        RECT 192.380 995.700 197.940 996.000 ;
        RECT 199.100 995.700 204.660 996.000 ;
        RECT 205.820 995.700 211.380 996.000 ;
        RECT 212.540 995.700 218.100 996.000 ;
        RECT 219.260 995.700 224.820 996.000 ;
        RECT 225.980 995.700 231.540 996.000 ;
        RECT 232.700 995.700 238.260 996.000 ;
        RECT 239.420 995.700 244.980 996.000 ;
        RECT 246.140 995.700 251.700 996.000 ;
        RECT 252.860 995.700 258.420 996.000 ;
        RECT 259.580 995.700 265.140 996.000 ;
        RECT 266.300 995.700 271.860 996.000 ;
        RECT 273.020 995.700 275.220 996.000 ;
        RECT 276.380 995.700 281.940 996.000 ;
        RECT 283.100 995.700 288.660 996.000 ;
        RECT 289.820 995.700 295.380 996.000 ;
        RECT 296.540 995.700 302.100 996.000 ;
        RECT 303.260 995.700 308.820 996.000 ;
        RECT 309.980 995.700 315.540 996.000 ;
        RECT 316.700 995.700 322.260 996.000 ;
        RECT 323.420 995.700 328.980 996.000 ;
        RECT 330.140 995.700 335.700 996.000 ;
        RECT 336.860 995.700 342.420 996.000 ;
        RECT 343.580 995.700 349.140 996.000 ;
        RECT 350.300 995.700 355.860 996.000 ;
        RECT 357.020 995.700 362.580 996.000 ;
        RECT 363.740 995.700 369.300 996.000 ;
        RECT 370.460 995.700 376.020 996.000 ;
        RECT 377.180 995.700 382.740 996.000 ;
        RECT 383.900 995.700 389.460 996.000 ;
        RECT 390.620 995.700 396.180 996.000 ;
        RECT 397.340 995.700 402.900 996.000 ;
        RECT 404.060 995.700 409.620 996.000 ;
        RECT 410.780 995.700 416.340 996.000 ;
        RECT 417.500 995.700 423.060 996.000 ;
        RECT 424.220 995.700 429.780 996.000 ;
        RECT 430.940 995.700 436.500 996.000 ;
        RECT 437.660 995.700 443.220 996.000 ;
        RECT 444.380 995.700 449.940 996.000 ;
        RECT 451.100 995.700 453.300 996.000 ;
        RECT 454.460 995.700 460.020 996.000 ;
        RECT 461.180 995.700 466.740 996.000 ;
        RECT 467.900 995.700 473.460 996.000 ;
        RECT 474.620 995.700 480.180 996.000 ;
        RECT 481.340 995.700 486.900 996.000 ;
        RECT 488.060 995.700 493.620 996.000 ;
        RECT 494.780 995.700 500.340 996.000 ;
        RECT 501.500 995.700 507.060 996.000 ;
        RECT 508.220 995.700 513.780 996.000 ;
        RECT 514.940 995.700 520.500 996.000 ;
        RECT 521.660 995.700 527.220 996.000 ;
        RECT 528.380 995.700 533.940 996.000 ;
        RECT 535.100 995.700 540.660 996.000 ;
        RECT 541.820 995.700 547.380 996.000 ;
        RECT 548.540 995.700 554.100 996.000 ;
        RECT 555.260 995.700 560.820 996.000 ;
        RECT 561.980 995.700 567.540 996.000 ;
        RECT 568.700 995.700 574.260 996.000 ;
        RECT 575.420 995.700 580.980 996.000 ;
        RECT 582.140 995.700 587.700 996.000 ;
        RECT 588.860 995.700 594.420 996.000 ;
        RECT 595.580 995.700 601.140 996.000 ;
        RECT 602.300 995.700 607.860 996.000 ;
        RECT 609.020 995.700 614.580 996.000 ;
        RECT 615.740 995.700 621.300 996.000 ;
        RECT 622.460 995.700 628.020 996.000 ;
        RECT 629.180 995.700 634.740 996.000 ;
        RECT 635.900 995.700 638.100 996.000 ;
        RECT 639.260 995.700 644.820 996.000 ;
        RECT 645.980 995.700 651.540 996.000 ;
        RECT 652.700 995.700 658.260 996.000 ;
        RECT 659.420 995.700 664.980 996.000 ;
        RECT 666.140 995.700 671.700 996.000 ;
        RECT 672.860 995.700 678.420 996.000 ;
        RECT 679.580 995.700 685.140 996.000 ;
        RECT 686.300 995.700 691.860 996.000 ;
        RECT 693.020 995.700 698.580 996.000 ;
        RECT 699.740 995.700 705.300 996.000 ;
        RECT 706.460 995.700 712.020 996.000 ;
        RECT 713.180 995.700 718.740 996.000 ;
        RECT 719.900 995.700 725.460 996.000 ;
        RECT 726.620 995.700 732.180 996.000 ;
        RECT 733.340 995.700 738.900 996.000 ;
        RECT 740.060 995.700 745.620 996.000 ;
        RECT 746.780 995.700 752.340 996.000 ;
        RECT 753.500 995.700 759.060 996.000 ;
        RECT 760.220 995.700 765.780 996.000 ;
        RECT 766.940 995.700 772.500 996.000 ;
        RECT 773.660 995.700 779.220 996.000 ;
        RECT 780.380 995.700 785.940 996.000 ;
        RECT 787.100 995.700 792.660 996.000 ;
        RECT 793.820 995.700 799.380 996.000 ;
        RECT 800.540 995.700 806.100 996.000 ;
        RECT 807.260 995.700 812.820 996.000 ;
        RECT 813.980 995.700 816.180 996.000 ;
        RECT 817.340 995.700 822.900 996.000 ;
        RECT 824.060 995.700 829.620 996.000 ;
        RECT 830.780 995.700 836.340 996.000 ;
        RECT 837.500 995.700 843.060 996.000 ;
        RECT 844.220 995.700 849.780 996.000 ;
        RECT 850.940 995.700 856.500 996.000 ;
        RECT 857.660 995.700 863.220 996.000 ;
        RECT 864.380 995.700 869.940 996.000 ;
        RECT 871.100 995.700 876.660 996.000 ;
        RECT 877.820 995.700 883.380 996.000 ;
        RECT 884.540 995.700 890.100 996.000 ;
        RECT 891.260 995.700 896.820 996.000 ;
        RECT 897.980 995.700 903.540 996.000 ;
        RECT 904.700 995.700 910.260 996.000 ;
        RECT 911.420 995.700 916.980 996.000 ;
        RECT 918.140 995.700 923.700 996.000 ;
        RECT 924.860 995.700 930.420 996.000 ;
        RECT 931.580 995.700 937.140 996.000 ;
        RECT 938.300 995.700 943.860 996.000 ;
        RECT 945.020 995.700 950.580 996.000 ;
        RECT 951.740 995.700 957.300 996.000 ;
        RECT 958.460 995.700 964.020 996.000 ;
        RECT 965.180 995.700 970.740 996.000 ;
        RECT 971.900 995.700 977.460 996.000 ;
        RECT 978.620 995.700 984.180 996.000 ;
        RECT 985.340 995.700 990.900 996.000 ;
        RECT 0.140 4.300 991.620 995.700 ;
        RECT 0.860 0.700 3.060 4.300 ;
        RECT 4.220 0.700 9.780 4.300 ;
        RECT 10.940 0.700 16.500 4.300 ;
        RECT 17.660 0.700 23.220 4.300 ;
        RECT 24.380 0.700 29.940 4.300 ;
        RECT 31.100 0.700 36.660 4.300 ;
        RECT 37.820 0.700 43.380 4.300 ;
        RECT 44.540 0.700 50.100 4.300 ;
        RECT 51.260 0.700 56.820 4.300 ;
        RECT 57.980 0.700 63.540 4.300 ;
        RECT 64.700 0.700 70.260 4.300 ;
        RECT 71.420 0.700 76.980 4.300 ;
        RECT 78.140 0.700 83.700 4.300 ;
        RECT 84.860 0.700 90.420 4.300 ;
        RECT 91.580 0.700 97.140 4.300 ;
        RECT 98.300 0.700 103.860 4.300 ;
        RECT 105.020 0.700 110.580 4.300 ;
        RECT 111.740 0.700 117.300 4.300 ;
        RECT 118.460 0.700 124.020 4.300 ;
        RECT 125.180 0.700 130.740 4.300 ;
        RECT 131.900 0.700 137.460 4.300 ;
        RECT 138.620 0.700 144.180 4.300 ;
        RECT 145.340 0.700 150.900 4.300 ;
        RECT 152.060 0.700 157.620 4.300 ;
        RECT 158.780 0.700 164.340 4.300 ;
        RECT 165.500 0.700 171.060 4.300 ;
        RECT 172.220 0.700 177.780 4.300 ;
        RECT 178.940 0.700 181.140 4.300 ;
        RECT 182.300 0.700 187.860 4.300 ;
        RECT 189.020 0.700 194.580 4.300 ;
        RECT 195.740 0.700 201.300 4.300 ;
        RECT 202.460 0.700 208.020 4.300 ;
        RECT 209.180 0.700 214.740 4.300 ;
        RECT 215.900 0.700 221.460 4.300 ;
        RECT 222.620 0.700 228.180 4.300 ;
        RECT 229.340 0.700 234.900 4.300 ;
        RECT 236.060 0.700 241.620 4.300 ;
        RECT 242.780 0.700 248.340 4.300 ;
        RECT 249.500 0.700 255.060 4.300 ;
        RECT 256.220 0.700 261.780 4.300 ;
        RECT 262.940 0.700 268.500 4.300 ;
        RECT 269.660 0.700 275.220 4.300 ;
        RECT 276.380 0.700 281.940 4.300 ;
        RECT 283.100 0.700 288.660 4.300 ;
        RECT 289.820 0.700 295.380 4.300 ;
        RECT 296.540 0.700 302.100 4.300 ;
        RECT 303.260 0.700 308.820 4.300 ;
        RECT 309.980 0.700 315.540 4.300 ;
        RECT 316.700 0.700 322.260 4.300 ;
        RECT 323.420 0.700 328.980 4.300 ;
        RECT 330.140 0.700 335.700 4.300 ;
        RECT 336.860 0.700 342.420 4.300 ;
        RECT 343.580 0.700 349.140 4.300 ;
        RECT 350.300 0.700 355.860 4.300 ;
        RECT 357.020 0.700 362.580 4.300 ;
        RECT 363.740 0.700 365.940 4.300 ;
        RECT 367.100 0.700 372.660 4.300 ;
        RECT 373.820 0.700 379.380 4.300 ;
        RECT 380.540 0.700 386.100 4.300 ;
        RECT 387.260 0.700 392.820 4.300 ;
        RECT 393.980 0.700 399.540 4.300 ;
        RECT 400.700 0.700 406.260 4.300 ;
        RECT 407.420 0.700 412.980 4.300 ;
        RECT 414.140 0.700 419.700 4.300 ;
        RECT 420.860 0.700 426.420 4.300 ;
        RECT 427.580 0.700 433.140 4.300 ;
        RECT 434.300 0.700 439.860 4.300 ;
        RECT 441.020 0.700 446.580 4.300 ;
        RECT 447.740 0.700 453.300 4.300 ;
        RECT 454.460 0.700 460.020 4.300 ;
        RECT 461.180 0.700 466.740 4.300 ;
        RECT 467.900 0.700 473.460 4.300 ;
        RECT 474.620 0.700 480.180 4.300 ;
        RECT 481.340 0.700 486.900 4.300 ;
        RECT 488.060 0.700 493.620 4.300 ;
        RECT 494.780 0.700 500.340 4.300 ;
        RECT 501.500 0.700 507.060 4.300 ;
        RECT 508.220 0.700 513.780 4.300 ;
        RECT 514.940 0.700 520.500 4.300 ;
        RECT 521.660 0.700 527.220 4.300 ;
        RECT 528.380 0.700 533.940 4.300 ;
        RECT 535.100 0.700 540.660 4.300 ;
        RECT 541.820 0.700 544.020 4.300 ;
        RECT 545.180 0.700 550.740 4.300 ;
        RECT 551.900 0.700 557.460 4.300 ;
        RECT 558.620 0.700 564.180 4.300 ;
        RECT 565.340 0.700 570.900 4.300 ;
        RECT 572.060 0.700 577.620 4.300 ;
        RECT 578.780 0.700 584.340 4.300 ;
        RECT 585.500 0.700 591.060 4.300 ;
        RECT 592.220 0.700 597.780 4.300 ;
        RECT 598.940 0.700 604.500 4.300 ;
        RECT 605.660 0.700 611.220 4.300 ;
        RECT 612.380 0.700 617.940 4.300 ;
        RECT 619.100 0.700 624.660 4.300 ;
        RECT 625.820 0.700 631.380 4.300 ;
        RECT 632.540 0.700 638.100 4.300 ;
        RECT 639.260 0.700 644.820 4.300 ;
        RECT 645.980 0.700 651.540 4.300 ;
        RECT 652.700 0.700 658.260 4.300 ;
        RECT 659.420 0.700 664.980 4.300 ;
        RECT 666.140 0.700 671.700 4.300 ;
        RECT 672.860 0.700 678.420 4.300 ;
        RECT 679.580 0.700 685.140 4.300 ;
        RECT 686.300 0.700 691.860 4.300 ;
        RECT 693.020 0.700 698.580 4.300 ;
        RECT 699.740 0.700 705.300 4.300 ;
        RECT 706.460 0.700 712.020 4.300 ;
        RECT 713.180 0.700 718.740 4.300 ;
        RECT 719.900 0.700 725.460 4.300 ;
        RECT 726.620 0.700 728.820 4.300 ;
        RECT 729.980 0.700 735.540 4.300 ;
        RECT 736.700 0.700 742.260 4.300 ;
        RECT 743.420 0.700 748.980 4.300 ;
        RECT 750.140 0.700 755.700 4.300 ;
        RECT 756.860 0.700 762.420 4.300 ;
        RECT 763.580 0.700 769.140 4.300 ;
        RECT 770.300 0.700 775.860 4.300 ;
        RECT 777.020 0.700 782.580 4.300 ;
        RECT 783.740 0.700 789.300 4.300 ;
        RECT 790.460 0.700 796.020 4.300 ;
        RECT 797.180 0.700 802.740 4.300 ;
        RECT 803.900 0.700 809.460 4.300 ;
        RECT 810.620 0.700 816.180 4.300 ;
        RECT 817.340 0.700 822.900 4.300 ;
        RECT 824.060 0.700 829.620 4.300 ;
        RECT 830.780 0.700 836.340 4.300 ;
        RECT 837.500 0.700 843.060 4.300 ;
        RECT 844.220 0.700 849.780 4.300 ;
        RECT 850.940 0.700 856.500 4.300 ;
        RECT 857.660 0.700 863.220 4.300 ;
        RECT 864.380 0.700 869.940 4.300 ;
        RECT 871.100 0.700 876.660 4.300 ;
        RECT 877.820 0.700 883.380 4.300 ;
        RECT 884.540 0.700 890.100 4.300 ;
        RECT 891.260 0.700 896.820 4.300 ;
        RECT 897.980 0.700 903.540 4.300 ;
        RECT 904.700 0.700 906.900 4.300 ;
        RECT 908.060 0.700 913.620 4.300 ;
        RECT 914.780 0.700 920.340 4.300 ;
        RECT 921.500 0.700 927.060 4.300 ;
        RECT 928.220 0.700 933.780 4.300 ;
        RECT 934.940 0.700 940.500 4.300 ;
        RECT 941.660 0.700 947.220 4.300 ;
        RECT 948.380 0.700 953.940 4.300 ;
        RECT 955.100 0.700 960.660 4.300 ;
        RECT 961.820 0.700 967.380 4.300 ;
        RECT 968.540 0.700 974.100 4.300 ;
        RECT 975.260 0.700 980.820 4.300 ;
        RECT 981.980 0.700 987.540 4.300 ;
        RECT 988.700 0.700 991.620 4.300 ;
        RECT 0.140 0.090 991.620 0.700 ;
      LAYER Metal3 ;
        RECT 0.090 990.900 995.700 991.620 ;
        RECT 0.090 988.700 996.000 990.900 ;
        RECT 0.090 987.540 0.700 988.700 ;
        RECT 4.300 987.540 996.000 988.700 ;
        RECT 0.090 985.340 996.000 987.540 ;
        RECT 0.090 984.180 995.700 985.340 ;
        RECT 0.090 981.980 996.000 984.180 ;
        RECT 0.090 980.820 0.700 981.980 ;
        RECT 4.300 980.820 996.000 981.980 ;
        RECT 0.090 978.620 996.000 980.820 ;
        RECT 0.090 977.460 995.700 978.620 ;
        RECT 0.090 975.260 996.000 977.460 ;
        RECT 0.090 974.100 0.700 975.260 ;
        RECT 4.300 974.100 996.000 975.260 ;
        RECT 0.090 971.900 996.000 974.100 ;
        RECT 0.090 970.740 995.700 971.900 ;
        RECT 0.090 968.540 996.000 970.740 ;
        RECT 0.090 967.380 0.700 968.540 ;
        RECT 4.300 967.380 996.000 968.540 ;
        RECT 0.090 965.180 996.000 967.380 ;
        RECT 0.090 964.020 995.700 965.180 ;
        RECT 0.090 961.820 996.000 964.020 ;
        RECT 0.090 960.660 0.700 961.820 ;
        RECT 4.300 960.660 996.000 961.820 ;
        RECT 0.090 958.460 996.000 960.660 ;
        RECT 0.090 957.300 995.700 958.460 ;
        RECT 0.090 955.100 996.000 957.300 ;
        RECT 0.090 953.940 0.700 955.100 ;
        RECT 4.300 953.940 996.000 955.100 ;
        RECT 0.090 951.740 996.000 953.940 ;
        RECT 0.090 950.580 995.700 951.740 ;
        RECT 0.090 948.380 996.000 950.580 ;
        RECT 0.090 947.220 0.700 948.380 ;
        RECT 4.300 947.220 996.000 948.380 ;
        RECT 0.090 945.020 996.000 947.220 ;
        RECT 0.090 943.860 995.700 945.020 ;
        RECT 0.090 941.660 996.000 943.860 ;
        RECT 0.090 940.500 0.700 941.660 ;
        RECT 4.300 940.500 996.000 941.660 ;
        RECT 0.090 938.300 996.000 940.500 ;
        RECT 0.090 937.140 995.700 938.300 ;
        RECT 0.090 934.940 996.000 937.140 ;
        RECT 0.090 933.780 0.700 934.940 ;
        RECT 4.300 933.780 996.000 934.940 ;
        RECT 0.090 931.580 996.000 933.780 ;
        RECT 0.090 930.420 995.700 931.580 ;
        RECT 0.090 928.220 996.000 930.420 ;
        RECT 0.090 927.060 0.700 928.220 ;
        RECT 4.300 927.060 996.000 928.220 ;
        RECT 0.090 924.860 996.000 927.060 ;
        RECT 0.090 923.700 995.700 924.860 ;
        RECT 0.090 921.500 996.000 923.700 ;
        RECT 0.090 920.340 0.700 921.500 ;
        RECT 4.300 920.340 996.000 921.500 ;
        RECT 0.090 918.140 996.000 920.340 ;
        RECT 0.090 916.980 995.700 918.140 ;
        RECT 0.090 914.780 996.000 916.980 ;
        RECT 0.090 913.620 0.700 914.780 ;
        RECT 4.300 913.620 996.000 914.780 ;
        RECT 0.090 911.420 996.000 913.620 ;
        RECT 0.090 910.260 995.700 911.420 ;
        RECT 0.090 908.060 996.000 910.260 ;
        RECT 0.090 906.900 0.700 908.060 ;
        RECT 4.300 906.900 996.000 908.060 ;
        RECT 0.090 904.700 996.000 906.900 ;
        RECT 0.090 903.540 0.700 904.700 ;
        RECT 4.300 903.540 995.700 904.700 ;
        RECT 0.090 897.980 996.000 903.540 ;
        RECT 0.090 896.820 0.700 897.980 ;
        RECT 4.300 896.820 995.700 897.980 ;
        RECT 0.090 891.260 996.000 896.820 ;
        RECT 0.090 890.100 0.700 891.260 ;
        RECT 4.300 890.100 995.700 891.260 ;
        RECT 0.090 884.540 996.000 890.100 ;
        RECT 0.090 883.380 0.700 884.540 ;
        RECT 4.300 883.380 995.700 884.540 ;
        RECT 0.090 877.820 996.000 883.380 ;
        RECT 0.090 876.660 0.700 877.820 ;
        RECT 4.300 876.660 995.700 877.820 ;
        RECT 0.090 871.100 996.000 876.660 ;
        RECT 0.090 869.940 0.700 871.100 ;
        RECT 4.300 869.940 995.700 871.100 ;
        RECT 0.090 864.380 996.000 869.940 ;
        RECT 0.090 863.220 0.700 864.380 ;
        RECT 4.300 863.220 995.700 864.380 ;
        RECT 0.090 857.660 996.000 863.220 ;
        RECT 0.090 856.500 0.700 857.660 ;
        RECT 4.300 856.500 995.700 857.660 ;
        RECT 0.090 850.940 996.000 856.500 ;
        RECT 0.090 849.780 0.700 850.940 ;
        RECT 4.300 849.780 995.700 850.940 ;
        RECT 0.090 844.220 996.000 849.780 ;
        RECT 0.090 843.060 0.700 844.220 ;
        RECT 4.300 843.060 995.700 844.220 ;
        RECT 0.090 837.500 996.000 843.060 ;
        RECT 0.090 836.340 0.700 837.500 ;
        RECT 4.300 836.340 995.700 837.500 ;
        RECT 0.090 830.780 996.000 836.340 ;
        RECT 0.090 829.620 0.700 830.780 ;
        RECT 4.300 829.620 995.700 830.780 ;
        RECT 0.090 824.060 996.000 829.620 ;
        RECT 0.090 822.900 0.700 824.060 ;
        RECT 4.300 822.900 995.700 824.060 ;
        RECT 0.090 817.340 996.000 822.900 ;
        RECT 0.090 816.180 0.700 817.340 ;
        RECT 4.300 816.180 995.700 817.340 ;
        RECT 0.090 813.980 996.000 816.180 ;
        RECT 0.090 812.820 995.700 813.980 ;
        RECT 0.090 810.620 996.000 812.820 ;
        RECT 0.090 809.460 0.700 810.620 ;
        RECT 4.300 809.460 996.000 810.620 ;
        RECT 0.090 807.260 996.000 809.460 ;
        RECT 0.090 806.100 995.700 807.260 ;
        RECT 0.090 803.900 996.000 806.100 ;
        RECT 0.090 802.740 0.700 803.900 ;
        RECT 4.300 802.740 996.000 803.900 ;
        RECT 0.090 800.540 996.000 802.740 ;
        RECT 0.090 799.380 995.700 800.540 ;
        RECT 0.090 797.180 996.000 799.380 ;
        RECT 0.090 796.020 0.700 797.180 ;
        RECT 4.300 796.020 996.000 797.180 ;
        RECT 0.090 793.820 996.000 796.020 ;
        RECT 0.090 792.660 995.700 793.820 ;
        RECT 0.090 790.460 996.000 792.660 ;
        RECT 0.090 789.300 0.700 790.460 ;
        RECT 4.300 789.300 996.000 790.460 ;
        RECT 0.090 787.100 996.000 789.300 ;
        RECT 0.090 785.940 995.700 787.100 ;
        RECT 0.090 783.740 996.000 785.940 ;
        RECT 0.090 782.580 0.700 783.740 ;
        RECT 4.300 782.580 996.000 783.740 ;
        RECT 0.090 780.380 996.000 782.580 ;
        RECT 0.090 779.220 995.700 780.380 ;
        RECT 0.090 777.020 996.000 779.220 ;
        RECT 0.090 775.860 0.700 777.020 ;
        RECT 4.300 775.860 996.000 777.020 ;
        RECT 0.090 773.660 996.000 775.860 ;
        RECT 0.090 772.500 995.700 773.660 ;
        RECT 0.090 770.300 996.000 772.500 ;
        RECT 0.090 769.140 0.700 770.300 ;
        RECT 4.300 769.140 996.000 770.300 ;
        RECT 0.090 766.940 996.000 769.140 ;
        RECT 0.090 765.780 995.700 766.940 ;
        RECT 0.090 763.580 996.000 765.780 ;
        RECT 0.090 762.420 0.700 763.580 ;
        RECT 4.300 762.420 996.000 763.580 ;
        RECT 0.090 760.220 996.000 762.420 ;
        RECT 0.090 759.060 995.700 760.220 ;
        RECT 0.090 756.860 996.000 759.060 ;
        RECT 0.090 755.700 0.700 756.860 ;
        RECT 4.300 755.700 996.000 756.860 ;
        RECT 0.090 753.500 996.000 755.700 ;
        RECT 0.090 752.340 995.700 753.500 ;
        RECT 0.090 750.140 996.000 752.340 ;
        RECT 0.090 748.980 0.700 750.140 ;
        RECT 4.300 748.980 996.000 750.140 ;
        RECT 0.090 746.780 996.000 748.980 ;
        RECT 0.090 745.620 995.700 746.780 ;
        RECT 0.090 743.420 996.000 745.620 ;
        RECT 0.090 742.260 0.700 743.420 ;
        RECT 4.300 742.260 996.000 743.420 ;
        RECT 0.090 740.060 996.000 742.260 ;
        RECT 0.090 738.900 995.700 740.060 ;
        RECT 0.090 736.700 996.000 738.900 ;
        RECT 0.090 735.540 0.700 736.700 ;
        RECT 4.300 735.540 996.000 736.700 ;
        RECT 0.090 733.340 996.000 735.540 ;
        RECT 0.090 732.180 995.700 733.340 ;
        RECT 0.090 729.980 996.000 732.180 ;
        RECT 0.090 728.820 0.700 729.980 ;
        RECT 4.300 728.820 996.000 729.980 ;
        RECT 0.090 726.620 996.000 728.820 ;
        RECT 0.090 725.460 0.700 726.620 ;
        RECT 4.300 725.460 995.700 726.620 ;
        RECT 0.090 719.900 996.000 725.460 ;
        RECT 0.090 718.740 0.700 719.900 ;
        RECT 4.300 718.740 995.700 719.900 ;
        RECT 0.090 713.180 996.000 718.740 ;
        RECT 0.090 712.020 0.700 713.180 ;
        RECT 4.300 712.020 995.700 713.180 ;
        RECT 0.090 706.460 996.000 712.020 ;
        RECT 0.090 705.300 0.700 706.460 ;
        RECT 4.300 705.300 995.700 706.460 ;
        RECT 0.090 699.740 996.000 705.300 ;
        RECT 0.090 698.580 0.700 699.740 ;
        RECT 4.300 698.580 995.700 699.740 ;
        RECT 0.090 693.020 996.000 698.580 ;
        RECT 0.090 691.860 0.700 693.020 ;
        RECT 4.300 691.860 995.700 693.020 ;
        RECT 0.090 686.300 996.000 691.860 ;
        RECT 0.090 685.140 0.700 686.300 ;
        RECT 4.300 685.140 995.700 686.300 ;
        RECT 0.090 679.580 996.000 685.140 ;
        RECT 0.090 678.420 0.700 679.580 ;
        RECT 4.300 678.420 995.700 679.580 ;
        RECT 0.090 672.860 996.000 678.420 ;
        RECT 0.090 671.700 0.700 672.860 ;
        RECT 4.300 671.700 995.700 672.860 ;
        RECT 0.090 666.140 996.000 671.700 ;
        RECT 0.090 664.980 0.700 666.140 ;
        RECT 4.300 664.980 995.700 666.140 ;
        RECT 0.090 659.420 996.000 664.980 ;
        RECT 0.090 658.260 0.700 659.420 ;
        RECT 4.300 658.260 995.700 659.420 ;
        RECT 0.090 652.700 996.000 658.260 ;
        RECT 0.090 651.540 0.700 652.700 ;
        RECT 4.300 651.540 995.700 652.700 ;
        RECT 0.090 645.980 996.000 651.540 ;
        RECT 0.090 644.820 0.700 645.980 ;
        RECT 4.300 644.820 995.700 645.980 ;
        RECT 0.090 639.260 996.000 644.820 ;
        RECT 0.090 638.100 0.700 639.260 ;
        RECT 4.300 638.100 995.700 639.260 ;
        RECT 0.090 635.900 996.000 638.100 ;
        RECT 0.090 634.740 995.700 635.900 ;
        RECT 0.090 632.540 996.000 634.740 ;
        RECT 0.090 631.380 0.700 632.540 ;
        RECT 4.300 631.380 996.000 632.540 ;
        RECT 0.090 629.180 996.000 631.380 ;
        RECT 0.090 628.020 995.700 629.180 ;
        RECT 0.090 625.820 996.000 628.020 ;
        RECT 0.090 624.660 0.700 625.820 ;
        RECT 4.300 624.660 996.000 625.820 ;
        RECT 0.090 622.460 996.000 624.660 ;
        RECT 0.090 621.300 995.700 622.460 ;
        RECT 0.090 619.100 996.000 621.300 ;
        RECT 0.090 617.940 0.700 619.100 ;
        RECT 4.300 617.940 996.000 619.100 ;
        RECT 0.090 615.740 996.000 617.940 ;
        RECT 0.090 614.580 995.700 615.740 ;
        RECT 0.090 612.380 996.000 614.580 ;
        RECT 0.090 611.220 0.700 612.380 ;
        RECT 4.300 611.220 996.000 612.380 ;
        RECT 0.090 609.020 996.000 611.220 ;
        RECT 0.090 607.860 995.700 609.020 ;
        RECT 0.090 605.660 996.000 607.860 ;
        RECT 0.090 604.500 0.700 605.660 ;
        RECT 4.300 604.500 996.000 605.660 ;
        RECT 0.090 602.300 996.000 604.500 ;
        RECT 0.090 601.140 995.700 602.300 ;
        RECT 0.090 598.940 996.000 601.140 ;
        RECT 0.090 597.780 0.700 598.940 ;
        RECT 4.300 597.780 996.000 598.940 ;
        RECT 0.090 595.580 996.000 597.780 ;
        RECT 0.090 594.420 995.700 595.580 ;
        RECT 0.090 592.220 996.000 594.420 ;
        RECT 0.090 591.060 0.700 592.220 ;
        RECT 4.300 591.060 996.000 592.220 ;
        RECT 0.090 588.860 996.000 591.060 ;
        RECT 0.090 587.700 995.700 588.860 ;
        RECT 0.090 585.500 996.000 587.700 ;
        RECT 0.090 584.340 0.700 585.500 ;
        RECT 4.300 584.340 996.000 585.500 ;
        RECT 0.090 582.140 996.000 584.340 ;
        RECT 0.090 580.980 995.700 582.140 ;
        RECT 0.090 578.780 996.000 580.980 ;
        RECT 0.090 577.620 0.700 578.780 ;
        RECT 4.300 577.620 996.000 578.780 ;
        RECT 0.090 575.420 996.000 577.620 ;
        RECT 0.090 574.260 995.700 575.420 ;
        RECT 0.090 572.060 996.000 574.260 ;
        RECT 0.090 570.900 0.700 572.060 ;
        RECT 4.300 570.900 996.000 572.060 ;
        RECT 0.090 568.700 996.000 570.900 ;
        RECT 0.090 567.540 995.700 568.700 ;
        RECT 0.090 565.340 996.000 567.540 ;
        RECT 0.090 564.180 0.700 565.340 ;
        RECT 4.300 564.180 996.000 565.340 ;
        RECT 0.090 561.980 996.000 564.180 ;
        RECT 0.090 560.820 995.700 561.980 ;
        RECT 0.090 558.620 996.000 560.820 ;
        RECT 0.090 557.460 0.700 558.620 ;
        RECT 4.300 557.460 996.000 558.620 ;
        RECT 0.090 555.260 996.000 557.460 ;
        RECT 0.090 554.100 995.700 555.260 ;
        RECT 0.090 551.900 996.000 554.100 ;
        RECT 0.090 550.740 0.700 551.900 ;
        RECT 4.300 550.740 996.000 551.900 ;
        RECT 0.090 548.540 996.000 550.740 ;
        RECT 0.090 547.380 995.700 548.540 ;
        RECT 0.090 545.180 996.000 547.380 ;
        RECT 0.090 544.020 0.700 545.180 ;
        RECT 4.300 544.020 996.000 545.180 ;
        RECT 0.090 541.820 996.000 544.020 ;
        RECT 0.090 540.660 0.700 541.820 ;
        RECT 4.300 540.660 995.700 541.820 ;
        RECT 0.090 535.100 996.000 540.660 ;
        RECT 0.090 533.940 0.700 535.100 ;
        RECT 4.300 533.940 995.700 535.100 ;
        RECT 0.090 528.380 996.000 533.940 ;
        RECT 0.090 527.220 0.700 528.380 ;
        RECT 4.300 527.220 995.700 528.380 ;
        RECT 0.090 521.660 996.000 527.220 ;
        RECT 0.090 520.500 0.700 521.660 ;
        RECT 4.300 520.500 995.700 521.660 ;
        RECT 0.090 514.940 996.000 520.500 ;
        RECT 0.090 513.780 0.700 514.940 ;
        RECT 4.300 513.780 995.700 514.940 ;
        RECT 0.090 508.220 996.000 513.780 ;
        RECT 0.090 507.060 0.700 508.220 ;
        RECT 4.300 507.060 995.700 508.220 ;
        RECT 0.090 501.500 996.000 507.060 ;
        RECT 0.090 500.340 0.700 501.500 ;
        RECT 4.300 500.340 995.700 501.500 ;
        RECT 0.090 494.780 996.000 500.340 ;
        RECT 0.090 493.620 0.700 494.780 ;
        RECT 4.300 493.620 995.700 494.780 ;
        RECT 0.090 488.060 996.000 493.620 ;
        RECT 0.090 486.900 0.700 488.060 ;
        RECT 4.300 486.900 995.700 488.060 ;
        RECT 0.090 481.340 996.000 486.900 ;
        RECT 0.090 480.180 0.700 481.340 ;
        RECT 4.300 480.180 995.700 481.340 ;
        RECT 0.090 474.620 996.000 480.180 ;
        RECT 0.090 473.460 0.700 474.620 ;
        RECT 4.300 473.460 995.700 474.620 ;
        RECT 0.090 467.900 996.000 473.460 ;
        RECT 0.090 466.740 0.700 467.900 ;
        RECT 4.300 466.740 995.700 467.900 ;
        RECT 0.090 461.180 996.000 466.740 ;
        RECT 0.090 460.020 0.700 461.180 ;
        RECT 4.300 460.020 995.700 461.180 ;
        RECT 0.090 454.460 996.000 460.020 ;
        RECT 0.090 453.300 0.700 454.460 ;
        RECT 4.300 453.300 995.700 454.460 ;
        RECT 0.090 451.100 996.000 453.300 ;
        RECT 0.090 449.940 995.700 451.100 ;
        RECT 0.090 447.740 996.000 449.940 ;
        RECT 0.090 446.580 0.700 447.740 ;
        RECT 4.300 446.580 996.000 447.740 ;
        RECT 0.090 444.380 996.000 446.580 ;
        RECT 0.090 443.220 995.700 444.380 ;
        RECT 0.090 441.020 996.000 443.220 ;
        RECT 0.090 439.860 0.700 441.020 ;
        RECT 4.300 439.860 996.000 441.020 ;
        RECT 0.090 437.660 996.000 439.860 ;
        RECT 0.090 436.500 995.700 437.660 ;
        RECT 0.090 434.300 996.000 436.500 ;
        RECT 0.090 433.140 0.700 434.300 ;
        RECT 4.300 433.140 996.000 434.300 ;
        RECT 0.090 430.940 996.000 433.140 ;
        RECT 0.090 429.780 995.700 430.940 ;
        RECT 0.090 427.580 996.000 429.780 ;
        RECT 0.090 426.420 0.700 427.580 ;
        RECT 4.300 426.420 996.000 427.580 ;
        RECT 0.090 424.220 996.000 426.420 ;
        RECT 0.090 423.060 995.700 424.220 ;
        RECT 0.090 420.860 996.000 423.060 ;
        RECT 0.090 419.700 0.700 420.860 ;
        RECT 4.300 419.700 996.000 420.860 ;
        RECT 0.090 417.500 996.000 419.700 ;
        RECT 0.090 416.340 995.700 417.500 ;
        RECT 0.090 414.140 996.000 416.340 ;
        RECT 0.090 412.980 0.700 414.140 ;
        RECT 4.300 412.980 996.000 414.140 ;
        RECT 0.090 410.780 996.000 412.980 ;
        RECT 0.090 409.620 995.700 410.780 ;
        RECT 0.090 407.420 996.000 409.620 ;
        RECT 0.090 406.260 0.700 407.420 ;
        RECT 4.300 406.260 996.000 407.420 ;
        RECT 0.090 404.060 996.000 406.260 ;
        RECT 0.090 402.900 995.700 404.060 ;
        RECT 0.090 400.700 996.000 402.900 ;
        RECT 0.090 399.540 0.700 400.700 ;
        RECT 4.300 399.540 996.000 400.700 ;
        RECT 0.090 397.340 996.000 399.540 ;
        RECT 0.090 396.180 995.700 397.340 ;
        RECT 0.090 393.980 996.000 396.180 ;
        RECT 0.090 392.820 0.700 393.980 ;
        RECT 4.300 392.820 996.000 393.980 ;
        RECT 0.090 390.620 996.000 392.820 ;
        RECT 0.090 389.460 995.700 390.620 ;
        RECT 0.090 387.260 996.000 389.460 ;
        RECT 0.090 386.100 0.700 387.260 ;
        RECT 4.300 386.100 996.000 387.260 ;
        RECT 0.090 383.900 996.000 386.100 ;
        RECT 0.090 382.740 995.700 383.900 ;
        RECT 0.090 380.540 996.000 382.740 ;
        RECT 0.090 379.380 0.700 380.540 ;
        RECT 4.300 379.380 996.000 380.540 ;
        RECT 0.090 377.180 996.000 379.380 ;
        RECT 0.090 376.020 995.700 377.180 ;
        RECT 0.090 373.820 996.000 376.020 ;
        RECT 0.090 372.660 0.700 373.820 ;
        RECT 4.300 372.660 996.000 373.820 ;
        RECT 0.090 370.460 996.000 372.660 ;
        RECT 0.090 369.300 995.700 370.460 ;
        RECT 0.090 367.100 996.000 369.300 ;
        RECT 0.090 365.940 0.700 367.100 ;
        RECT 4.300 365.940 996.000 367.100 ;
        RECT 0.090 363.740 996.000 365.940 ;
        RECT 0.090 362.580 0.700 363.740 ;
        RECT 4.300 362.580 995.700 363.740 ;
        RECT 0.090 357.020 996.000 362.580 ;
        RECT 0.090 355.860 0.700 357.020 ;
        RECT 4.300 355.860 995.700 357.020 ;
        RECT 0.090 350.300 996.000 355.860 ;
        RECT 0.090 349.140 0.700 350.300 ;
        RECT 4.300 349.140 995.700 350.300 ;
        RECT 0.090 343.580 996.000 349.140 ;
        RECT 0.090 342.420 0.700 343.580 ;
        RECT 4.300 342.420 995.700 343.580 ;
        RECT 0.090 336.860 996.000 342.420 ;
        RECT 0.090 335.700 0.700 336.860 ;
        RECT 4.300 335.700 995.700 336.860 ;
        RECT 0.090 330.140 996.000 335.700 ;
        RECT 0.090 328.980 0.700 330.140 ;
        RECT 4.300 328.980 995.700 330.140 ;
        RECT 0.090 323.420 996.000 328.980 ;
        RECT 0.090 322.260 0.700 323.420 ;
        RECT 4.300 322.260 995.700 323.420 ;
        RECT 0.090 316.700 996.000 322.260 ;
        RECT 0.090 315.540 0.700 316.700 ;
        RECT 4.300 315.540 995.700 316.700 ;
        RECT 0.090 309.980 996.000 315.540 ;
        RECT 0.090 308.820 0.700 309.980 ;
        RECT 4.300 308.820 995.700 309.980 ;
        RECT 0.090 303.260 996.000 308.820 ;
        RECT 0.090 302.100 0.700 303.260 ;
        RECT 4.300 302.100 995.700 303.260 ;
        RECT 0.090 296.540 996.000 302.100 ;
        RECT 0.090 295.380 0.700 296.540 ;
        RECT 4.300 295.380 995.700 296.540 ;
        RECT 0.090 289.820 996.000 295.380 ;
        RECT 0.090 288.660 0.700 289.820 ;
        RECT 4.300 288.660 995.700 289.820 ;
        RECT 0.090 283.100 996.000 288.660 ;
        RECT 0.090 281.940 0.700 283.100 ;
        RECT 4.300 281.940 995.700 283.100 ;
        RECT 0.090 276.380 996.000 281.940 ;
        RECT 0.090 275.220 0.700 276.380 ;
        RECT 4.300 275.220 995.700 276.380 ;
        RECT 0.090 273.020 996.000 275.220 ;
        RECT 0.090 271.860 995.700 273.020 ;
        RECT 0.090 269.660 996.000 271.860 ;
        RECT 0.090 268.500 0.700 269.660 ;
        RECT 4.300 268.500 996.000 269.660 ;
        RECT 0.090 266.300 996.000 268.500 ;
        RECT 0.090 265.140 995.700 266.300 ;
        RECT 0.090 262.940 996.000 265.140 ;
        RECT 0.090 261.780 0.700 262.940 ;
        RECT 4.300 261.780 996.000 262.940 ;
        RECT 0.090 259.580 996.000 261.780 ;
        RECT 0.090 258.420 995.700 259.580 ;
        RECT 0.090 256.220 996.000 258.420 ;
        RECT 0.090 255.060 0.700 256.220 ;
        RECT 4.300 255.060 996.000 256.220 ;
        RECT 0.090 252.860 996.000 255.060 ;
        RECT 0.090 251.700 995.700 252.860 ;
        RECT 0.090 249.500 996.000 251.700 ;
        RECT 0.090 248.340 0.700 249.500 ;
        RECT 4.300 248.340 996.000 249.500 ;
        RECT 0.090 246.140 996.000 248.340 ;
        RECT 0.090 244.980 995.700 246.140 ;
        RECT 0.090 242.780 996.000 244.980 ;
        RECT 0.090 241.620 0.700 242.780 ;
        RECT 4.300 241.620 996.000 242.780 ;
        RECT 0.090 239.420 996.000 241.620 ;
        RECT 0.090 238.260 995.700 239.420 ;
        RECT 0.090 236.060 996.000 238.260 ;
        RECT 0.090 234.900 0.700 236.060 ;
        RECT 4.300 234.900 996.000 236.060 ;
        RECT 0.090 232.700 996.000 234.900 ;
        RECT 0.090 231.540 995.700 232.700 ;
        RECT 0.090 229.340 996.000 231.540 ;
        RECT 0.090 228.180 0.700 229.340 ;
        RECT 4.300 228.180 996.000 229.340 ;
        RECT 0.090 225.980 996.000 228.180 ;
        RECT 0.090 224.820 995.700 225.980 ;
        RECT 0.090 222.620 996.000 224.820 ;
        RECT 0.090 221.460 0.700 222.620 ;
        RECT 4.300 221.460 996.000 222.620 ;
        RECT 0.090 219.260 996.000 221.460 ;
        RECT 0.090 218.100 995.700 219.260 ;
        RECT 0.090 215.900 996.000 218.100 ;
        RECT 0.090 214.740 0.700 215.900 ;
        RECT 4.300 214.740 996.000 215.900 ;
        RECT 0.090 212.540 996.000 214.740 ;
        RECT 0.090 211.380 995.700 212.540 ;
        RECT 0.090 209.180 996.000 211.380 ;
        RECT 0.090 208.020 0.700 209.180 ;
        RECT 4.300 208.020 996.000 209.180 ;
        RECT 0.090 205.820 996.000 208.020 ;
        RECT 0.090 204.660 995.700 205.820 ;
        RECT 0.090 202.460 996.000 204.660 ;
        RECT 0.090 201.300 0.700 202.460 ;
        RECT 4.300 201.300 996.000 202.460 ;
        RECT 0.090 199.100 996.000 201.300 ;
        RECT 0.090 197.940 995.700 199.100 ;
        RECT 0.090 195.740 996.000 197.940 ;
        RECT 0.090 194.580 0.700 195.740 ;
        RECT 4.300 194.580 996.000 195.740 ;
        RECT 0.090 192.380 996.000 194.580 ;
        RECT 0.090 191.220 995.700 192.380 ;
        RECT 0.090 189.020 996.000 191.220 ;
        RECT 0.090 187.860 0.700 189.020 ;
        RECT 4.300 187.860 996.000 189.020 ;
        RECT 0.090 185.660 996.000 187.860 ;
        RECT 0.090 184.500 995.700 185.660 ;
        RECT 0.090 182.300 996.000 184.500 ;
        RECT 0.090 181.140 0.700 182.300 ;
        RECT 4.300 181.140 996.000 182.300 ;
        RECT 0.090 178.940 996.000 181.140 ;
        RECT 0.090 177.780 0.700 178.940 ;
        RECT 4.300 177.780 995.700 178.940 ;
        RECT 0.090 172.220 996.000 177.780 ;
        RECT 0.090 171.060 0.700 172.220 ;
        RECT 4.300 171.060 995.700 172.220 ;
        RECT 0.090 165.500 996.000 171.060 ;
        RECT 0.090 164.340 0.700 165.500 ;
        RECT 4.300 164.340 995.700 165.500 ;
        RECT 0.090 158.780 996.000 164.340 ;
        RECT 0.090 157.620 0.700 158.780 ;
        RECT 4.300 157.620 995.700 158.780 ;
        RECT 0.090 152.060 996.000 157.620 ;
        RECT 0.090 150.900 0.700 152.060 ;
        RECT 4.300 150.900 995.700 152.060 ;
        RECT 0.090 145.340 996.000 150.900 ;
        RECT 0.090 144.180 0.700 145.340 ;
        RECT 4.300 144.180 995.700 145.340 ;
        RECT 0.090 138.620 996.000 144.180 ;
        RECT 0.090 137.460 0.700 138.620 ;
        RECT 4.300 137.460 995.700 138.620 ;
        RECT 0.090 131.900 996.000 137.460 ;
        RECT 0.090 130.740 0.700 131.900 ;
        RECT 4.300 130.740 995.700 131.900 ;
        RECT 0.090 125.180 996.000 130.740 ;
        RECT 0.090 124.020 0.700 125.180 ;
        RECT 4.300 124.020 995.700 125.180 ;
        RECT 0.090 118.460 996.000 124.020 ;
        RECT 0.090 117.300 0.700 118.460 ;
        RECT 4.300 117.300 995.700 118.460 ;
        RECT 0.090 111.740 996.000 117.300 ;
        RECT 0.090 110.580 0.700 111.740 ;
        RECT 4.300 110.580 995.700 111.740 ;
        RECT 0.090 105.020 996.000 110.580 ;
        RECT 0.090 103.860 0.700 105.020 ;
        RECT 4.300 103.860 995.700 105.020 ;
        RECT 0.090 98.300 996.000 103.860 ;
        RECT 0.090 97.140 0.700 98.300 ;
        RECT 4.300 97.140 995.700 98.300 ;
        RECT 0.090 91.580 996.000 97.140 ;
        RECT 0.090 90.420 0.700 91.580 ;
        RECT 4.300 90.420 995.700 91.580 ;
        RECT 0.090 88.220 996.000 90.420 ;
        RECT 0.090 87.060 995.700 88.220 ;
        RECT 0.090 84.860 996.000 87.060 ;
        RECT 0.090 83.700 0.700 84.860 ;
        RECT 4.300 83.700 996.000 84.860 ;
        RECT 0.090 81.500 996.000 83.700 ;
        RECT 0.090 80.340 995.700 81.500 ;
        RECT 0.090 78.140 996.000 80.340 ;
        RECT 0.090 76.980 0.700 78.140 ;
        RECT 4.300 76.980 996.000 78.140 ;
        RECT 0.090 74.780 996.000 76.980 ;
        RECT 0.090 73.620 995.700 74.780 ;
        RECT 0.090 71.420 996.000 73.620 ;
        RECT 0.090 70.260 0.700 71.420 ;
        RECT 4.300 70.260 996.000 71.420 ;
        RECT 0.090 68.060 996.000 70.260 ;
        RECT 0.090 66.900 995.700 68.060 ;
        RECT 0.090 64.700 996.000 66.900 ;
        RECT 0.090 63.540 0.700 64.700 ;
        RECT 4.300 63.540 996.000 64.700 ;
        RECT 0.090 61.340 996.000 63.540 ;
        RECT 0.090 60.180 995.700 61.340 ;
        RECT 0.090 57.980 996.000 60.180 ;
        RECT 0.090 56.820 0.700 57.980 ;
        RECT 4.300 56.820 996.000 57.980 ;
        RECT 0.090 54.620 996.000 56.820 ;
        RECT 0.090 53.460 995.700 54.620 ;
        RECT 0.090 51.260 996.000 53.460 ;
        RECT 0.090 50.100 0.700 51.260 ;
        RECT 4.300 50.100 996.000 51.260 ;
        RECT 0.090 47.900 996.000 50.100 ;
        RECT 0.090 46.740 995.700 47.900 ;
        RECT 0.090 44.540 996.000 46.740 ;
        RECT 0.090 43.380 0.700 44.540 ;
        RECT 4.300 43.380 996.000 44.540 ;
        RECT 0.090 41.180 996.000 43.380 ;
        RECT 0.090 40.020 995.700 41.180 ;
        RECT 0.090 37.820 996.000 40.020 ;
        RECT 0.090 36.660 0.700 37.820 ;
        RECT 4.300 36.660 996.000 37.820 ;
        RECT 0.090 34.460 996.000 36.660 ;
        RECT 0.090 33.300 995.700 34.460 ;
        RECT 0.090 31.100 996.000 33.300 ;
        RECT 0.090 29.940 0.700 31.100 ;
        RECT 4.300 29.940 996.000 31.100 ;
        RECT 0.090 27.740 996.000 29.940 ;
        RECT 0.090 26.580 995.700 27.740 ;
        RECT 0.090 24.380 996.000 26.580 ;
        RECT 0.090 23.220 0.700 24.380 ;
        RECT 4.300 23.220 996.000 24.380 ;
        RECT 0.090 21.020 996.000 23.220 ;
        RECT 0.090 19.860 995.700 21.020 ;
        RECT 0.090 17.660 996.000 19.860 ;
        RECT 0.090 16.500 0.700 17.660 ;
        RECT 4.300 16.500 996.000 17.660 ;
        RECT 0.090 14.300 996.000 16.500 ;
        RECT 0.090 13.140 995.700 14.300 ;
        RECT 0.090 10.940 996.000 13.140 ;
        RECT 0.090 9.780 0.700 10.940 ;
        RECT 4.300 9.780 996.000 10.940 ;
        RECT 0.090 7.580 996.000 9.780 ;
        RECT 0.090 6.420 995.700 7.580 ;
        RECT 0.090 4.220 996.000 6.420 ;
        RECT 0.090 3.060 0.700 4.220 ;
        RECT 4.300 3.060 996.000 4.220 ;
        RECT 0.090 0.860 996.000 3.060 ;
        RECT 0.090 0.140 995.700 0.860 ;
  END
END tiny_user_project
END LIBRARY

