magic
tech gf180mcuC
magscale 1 5
timestamp 1669733779
<< obsm1 >>
rect 672 855 99288 98422
<< metal2 >>
rect 0 99600 56 99900
rect 672 99600 728 99900
rect 1344 99600 1400 99900
rect 2016 99600 2072 99900
rect 2688 99600 2744 99900
rect 3360 99600 3416 99900
rect 4032 99600 4088 99900
rect 4704 99600 4760 99900
rect 5376 99600 5432 99900
rect 6048 99600 6104 99900
rect 6720 99600 6776 99900
rect 7392 99600 7448 99900
rect 8064 99600 8120 99900
rect 8736 99600 8792 99900
rect 9072 99600 9128 99900
rect 9744 99600 9800 99900
rect 10416 99600 10472 99900
rect 11088 99600 11144 99900
rect 11760 99600 11816 99900
rect 12432 99600 12488 99900
rect 13104 99600 13160 99900
rect 13776 99600 13832 99900
rect 14448 99600 14504 99900
rect 15120 99600 15176 99900
rect 15792 99600 15848 99900
rect 16464 99600 16520 99900
rect 17136 99600 17192 99900
rect 17808 99600 17864 99900
rect 18480 99600 18536 99900
rect 19152 99600 19208 99900
rect 19824 99600 19880 99900
rect 20496 99600 20552 99900
rect 21168 99600 21224 99900
rect 21840 99600 21896 99900
rect 22512 99600 22568 99900
rect 23184 99600 23240 99900
rect 23856 99600 23912 99900
rect 24528 99600 24584 99900
rect 25200 99600 25256 99900
rect 25872 99600 25928 99900
rect 26544 99600 26600 99900
rect 27216 99600 27272 99900
rect 27552 99600 27608 99900
rect 28224 99600 28280 99900
rect 28896 99600 28952 99900
rect 29568 99600 29624 99900
rect 30240 99600 30296 99900
rect 30912 99600 30968 99900
rect 31584 99600 31640 99900
rect 32256 99600 32312 99900
rect 32928 99600 32984 99900
rect 33600 99600 33656 99900
rect 34272 99600 34328 99900
rect 34944 99600 35000 99900
rect 35616 99600 35672 99900
rect 36288 99600 36344 99900
rect 36960 99600 37016 99900
rect 37632 99600 37688 99900
rect 38304 99600 38360 99900
rect 38976 99600 39032 99900
rect 39648 99600 39704 99900
rect 40320 99600 40376 99900
rect 40992 99600 41048 99900
rect 41664 99600 41720 99900
rect 42336 99600 42392 99900
rect 43008 99600 43064 99900
rect 43680 99600 43736 99900
rect 44352 99600 44408 99900
rect 45024 99600 45080 99900
rect 45360 99600 45416 99900
rect 46032 99600 46088 99900
rect 46704 99600 46760 99900
rect 47376 99600 47432 99900
rect 48048 99600 48104 99900
rect 48720 99600 48776 99900
rect 49392 99600 49448 99900
rect 50064 99600 50120 99900
rect 50736 99600 50792 99900
rect 51408 99600 51464 99900
rect 52080 99600 52136 99900
rect 52752 99600 52808 99900
rect 53424 99600 53480 99900
rect 54096 99600 54152 99900
rect 54768 99600 54824 99900
rect 55440 99600 55496 99900
rect 56112 99600 56168 99900
rect 56784 99600 56840 99900
rect 57456 99600 57512 99900
rect 58128 99600 58184 99900
rect 58800 99600 58856 99900
rect 59472 99600 59528 99900
rect 60144 99600 60200 99900
rect 60816 99600 60872 99900
rect 61488 99600 61544 99900
rect 62160 99600 62216 99900
rect 62832 99600 62888 99900
rect 63504 99600 63560 99900
rect 63840 99600 63896 99900
rect 64512 99600 64568 99900
rect 65184 99600 65240 99900
rect 65856 99600 65912 99900
rect 66528 99600 66584 99900
rect 67200 99600 67256 99900
rect 67872 99600 67928 99900
rect 68544 99600 68600 99900
rect 69216 99600 69272 99900
rect 69888 99600 69944 99900
rect 70560 99600 70616 99900
rect 71232 99600 71288 99900
rect 71904 99600 71960 99900
rect 72576 99600 72632 99900
rect 73248 99600 73304 99900
rect 73920 99600 73976 99900
rect 74592 99600 74648 99900
rect 75264 99600 75320 99900
rect 75936 99600 75992 99900
rect 76608 99600 76664 99900
rect 77280 99600 77336 99900
rect 77952 99600 78008 99900
rect 78624 99600 78680 99900
rect 79296 99600 79352 99900
rect 79968 99600 80024 99900
rect 80640 99600 80696 99900
rect 81312 99600 81368 99900
rect 81648 99600 81704 99900
rect 82320 99600 82376 99900
rect 82992 99600 83048 99900
rect 83664 99600 83720 99900
rect 84336 99600 84392 99900
rect 85008 99600 85064 99900
rect 85680 99600 85736 99900
rect 86352 99600 86408 99900
rect 87024 99600 87080 99900
rect 87696 99600 87752 99900
rect 88368 99600 88424 99900
rect 89040 99600 89096 99900
rect 89712 99600 89768 99900
rect 90384 99600 90440 99900
rect 91056 99600 91112 99900
rect 91728 99600 91784 99900
rect 92400 99600 92456 99900
rect 93072 99600 93128 99900
rect 93744 99600 93800 99900
rect 94416 99600 94472 99900
rect 95088 99600 95144 99900
rect 95760 99600 95816 99900
rect 96432 99600 96488 99900
rect 97104 99600 97160 99900
rect 97776 99600 97832 99900
rect 98448 99600 98504 99900
rect 99120 99600 99176 99900
rect 99792 99600 99848 99900
rect 0 100 56 400
rect 336 100 392 400
rect 1008 100 1064 400
rect 1680 100 1736 400
rect 2352 100 2408 400
rect 3024 100 3080 400
rect 3696 100 3752 400
rect 4368 100 4424 400
rect 5040 100 5096 400
rect 5712 100 5768 400
rect 6384 100 6440 400
rect 7056 100 7112 400
rect 7728 100 7784 400
rect 8400 100 8456 400
rect 9072 100 9128 400
rect 9744 100 9800 400
rect 10416 100 10472 400
rect 11088 100 11144 400
rect 11760 100 11816 400
rect 12432 100 12488 400
rect 13104 100 13160 400
rect 13776 100 13832 400
rect 14448 100 14504 400
rect 15120 100 15176 400
rect 15792 100 15848 400
rect 16464 100 16520 400
rect 17136 100 17192 400
rect 17808 100 17864 400
rect 18144 100 18200 400
rect 18816 100 18872 400
rect 19488 100 19544 400
rect 20160 100 20216 400
rect 20832 100 20888 400
rect 21504 100 21560 400
rect 22176 100 22232 400
rect 22848 100 22904 400
rect 23520 100 23576 400
rect 24192 100 24248 400
rect 24864 100 24920 400
rect 25536 100 25592 400
rect 26208 100 26264 400
rect 26880 100 26936 400
rect 27552 100 27608 400
rect 28224 100 28280 400
rect 28896 100 28952 400
rect 29568 100 29624 400
rect 30240 100 30296 400
rect 30912 100 30968 400
rect 31584 100 31640 400
rect 32256 100 32312 400
rect 32928 100 32984 400
rect 33600 100 33656 400
rect 34272 100 34328 400
rect 34944 100 35000 400
rect 35616 100 35672 400
rect 36288 100 36344 400
rect 36624 100 36680 400
rect 37296 100 37352 400
rect 37968 100 38024 400
rect 38640 100 38696 400
rect 39312 100 39368 400
rect 39984 100 40040 400
rect 40656 100 40712 400
rect 41328 100 41384 400
rect 42000 100 42056 400
rect 42672 100 42728 400
rect 43344 100 43400 400
rect 44016 100 44072 400
rect 44688 100 44744 400
rect 45360 100 45416 400
rect 46032 100 46088 400
rect 46704 100 46760 400
rect 47376 100 47432 400
rect 48048 100 48104 400
rect 48720 100 48776 400
rect 49392 100 49448 400
rect 50064 100 50120 400
rect 50736 100 50792 400
rect 51408 100 51464 400
rect 52080 100 52136 400
rect 52752 100 52808 400
rect 53424 100 53480 400
rect 54096 100 54152 400
rect 54432 100 54488 400
rect 55104 100 55160 400
rect 55776 100 55832 400
rect 56448 100 56504 400
rect 57120 100 57176 400
rect 57792 100 57848 400
rect 58464 100 58520 400
rect 59136 100 59192 400
rect 59808 100 59864 400
rect 60480 100 60536 400
rect 61152 100 61208 400
rect 61824 100 61880 400
rect 62496 100 62552 400
rect 63168 100 63224 400
rect 63840 100 63896 400
rect 64512 100 64568 400
rect 65184 100 65240 400
rect 65856 100 65912 400
rect 66528 100 66584 400
rect 67200 100 67256 400
rect 67872 100 67928 400
rect 68544 100 68600 400
rect 69216 100 69272 400
rect 69888 100 69944 400
rect 70560 100 70616 400
rect 71232 100 71288 400
rect 71904 100 71960 400
rect 72576 100 72632 400
rect 72912 100 72968 400
rect 73584 100 73640 400
rect 74256 100 74312 400
rect 74928 100 74984 400
rect 75600 100 75656 400
rect 76272 100 76328 400
rect 76944 100 77000 400
rect 77616 100 77672 400
rect 78288 100 78344 400
rect 78960 100 79016 400
rect 79632 100 79688 400
rect 80304 100 80360 400
rect 80976 100 81032 400
rect 81648 100 81704 400
rect 82320 100 82376 400
rect 82992 100 83048 400
rect 83664 100 83720 400
rect 84336 100 84392 400
rect 85008 100 85064 400
rect 85680 100 85736 400
rect 86352 100 86408 400
rect 87024 100 87080 400
rect 87696 100 87752 400
rect 88368 100 88424 400
rect 89040 100 89096 400
rect 89712 100 89768 400
rect 90384 100 90440 400
rect 90720 100 90776 400
rect 91392 100 91448 400
rect 92064 100 92120 400
rect 92736 100 92792 400
rect 93408 100 93464 400
rect 94080 100 94136 400
rect 94752 100 94808 400
rect 95424 100 95480 400
rect 96096 100 96152 400
rect 96768 100 96824 400
rect 97440 100 97496 400
rect 98112 100 98168 400
rect 98784 100 98840 400
rect 99456 100 99512 400
<< obsm2 >>
rect 86 99570 642 99600
rect 758 99570 1314 99600
rect 1430 99570 1986 99600
rect 2102 99570 2658 99600
rect 2774 99570 3330 99600
rect 3446 99570 4002 99600
rect 4118 99570 4674 99600
rect 4790 99570 5346 99600
rect 5462 99570 6018 99600
rect 6134 99570 6690 99600
rect 6806 99570 7362 99600
rect 7478 99570 8034 99600
rect 8150 99570 8706 99600
rect 8822 99570 9042 99600
rect 9158 99570 9714 99600
rect 9830 99570 10386 99600
rect 10502 99570 11058 99600
rect 11174 99570 11730 99600
rect 11846 99570 12402 99600
rect 12518 99570 13074 99600
rect 13190 99570 13746 99600
rect 13862 99570 14418 99600
rect 14534 99570 15090 99600
rect 15206 99570 15762 99600
rect 15878 99570 16434 99600
rect 16550 99570 17106 99600
rect 17222 99570 17778 99600
rect 17894 99570 18450 99600
rect 18566 99570 19122 99600
rect 19238 99570 19794 99600
rect 19910 99570 20466 99600
rect 20582 99570 21138 99600
rect 21254 99570 21810 99600
rect 21926 99570 22482 99600
rect 22598 99570 23154 99600
rect 23270 99570 23826 99600
rect 23942 99570 24498 99600
rect 24614 99570 25170 99600
rect 25286 99570 25842 99600
rect 25958 99570 26514 99600
rect 26630 99570 27186 99600
rect 27302 99570 27522 99600
rect 27638 99570 28194 99600
rect 28310 99570 28866 99600
rect 28982 99570 29538 99600
rect 29654 99570 30210 99600
rect 30326 99570 30882 99600
rect 30998 99570 31554 99600
rect 31670 99570 32226 99600
rect 32342 99570 32898 99600
rect 33014 99570 33570 99600
rect 33686 99570 34242 99600
rect 34358 99570 34914 99600
rect 35030 99570 35586 99600
rect 35702 99570 36258 99600
rect 36374 99570 36930 99600
rect 37046 99570 37602 99600
rect 37718 99570 38274 99600
rect 38390 99570 38946 99600
rect 39062 99570 39618 99600
rect 39734 99570 40290 99600
rect 40406 99570 40962 99600
rect 41078 99570 41634 99600
rect 41750 99570 42306 99600
rect 42422 99570 42978 99600
rect 43094 99570 43650 99600
rect 43766 99570 44322 99600
rect 44438 99570 44994 99600
rect 45110 99570 45330 99600
rect 45446 99570 46002 99600
rect 46118 99570 46674 99600
rect 46790 99570 47346 99600
rect 47462 99570 48018 99600
rect 48134 99570 48690 99600
rect 48806 99570 49362 99600
rect 49478 99570 50034 99600
rect 50150 99570 50706 99600
rect 50822 99570 51378 99600
rect 51494 99570 52050 99600
rect 52166 99570 52722 99600
rect 52838 99570 53394 99600
rect 53510 99570 54066 99600
rect 54182 99570 54738 99600
rect 54854 99570 55410 99600
rect 55526 99570 56082 99600
rect 56198 99570 56754 99600
rect 56870 99570 57426 99600
rect 57542 99570 58098 99600
rect 58214 99570 58770 99600
rect 58886 99570 59442 99600
rect 59558 99570 60114 99600
rect 60230 99570 60786 99600
rect 60902 99570 61458 99600
rect 61574 99570 62130 99600
rect 62246 99570 62802 99600
rect 62918 99570 63474 99600
rect 63590 99570 63810 99600
rect 63926 99570 64482 99600
rect 64598 99570 65154 99600
rect 65270 99570 65826 99600
rect 65942 99570 66498 99600
rect 66614 99570 67170 99600
rect 67286 99570 67842 99600
rect 67958 99570 68514 99600
rect 68630 99570 69186 99600
rect 69302 99570 69858 99600
rect 69974 99570 70530 99600
rect 70646 99570 71202 99600
rect 71318 99570 71874 99600
rect 71990 99570 72546 99600
rect 72662 99570 73218 99600
rect 73334 99570 73890 99600
rect 74006 99570 74562 99600
rect 74678 99570 75234 99600
rect 75350 99570 75906 99600
rect 76022 99570 76578 99600
rect 76694 99570 77250 99600
rect 77366 99570 77922 99600
rect 78038 99570 78594 99600
rect 78710 99570 79266 99600
rect 79382 99570 79938 99600
rect 80054 99570 80610 99600
rect 80726 99570 81282 99600
rect 81398 99570 81618 99600
rect 81734 99570 82290 99600
rect 82406 99570 82962 99600
rect 83078 99570 83634 99600
rect 83750 99570 84306 99600
rect 84422 99570 84978 99600
rect 85094 99570 85650 99600
rect 85766 99570 86322 99600
rect 86438 99570 86994 99600
rect 87110 99570 87666 99600
rect 87782 99570 88338 99600
rect 88454 99570 89010 99600
rect 89126 99570 89682 99600
rect 89798 99570 90354 99600
rect 90470 99570 91026 99600
rect 91142 99570 91698 99600
rect 91814 99570 92370 99600
rect 92486 99570 93042 99600
rect 93158 99570 93714 99600
rect 93830 99570 94386 99600
rect 94502 99570 95058 99600
rect 95174 99570 95730 99600
rect 95846 99570 96402 99600
rect 96518 99570 97074 99600
rect 97190 99570 97746 99600
rect 97862 99570 98418 99600
rect 98534 99570 99090 99600
rect 14 430 99162 99570
rect 86 70 306 430
rect 422 70 978 430
rect 1094 70 1650 430
rect 1766 70 2322 430
rect 2438 70 2994 430
rect 3110 70 3666 430
rect 3782 70 4338 430
rect 4454 70 5010 430
rect 5126 70 5682 430
rect 5798 70 6354 430
rect 6470 70 7026 430
rect 7142 70 7698 430
rect 7814 70 8370 430
rect 8486 70 9042 430
rect 9158 70 9714 430
rect 9830 70 10386 430
rect 10502 70 11058 430
rect 11174 70 11730 430
rect 11846 70 12402 430
rect 12518 70 13074 430
rect 13190 70 13746 430
rect 13862 70 14418 430
rect 14534 70 15090 430
rect 15206 70 15762 430
rect 15878 70 16434 430
rect 16550 70 17106 430
rect 17222 70 17778 430
rect 17894 70 18114 430
rect 18230 70 18786 430
rect 18902 70 19458 430
rect 19574 70 20130 430
rect 20246 70 20802 430
rect 20918 70 21474 430
rect 21590 70 22146 430
rect 22262 70 22818 430
rect 22934 70 23490 430
rect 23606 70 24162 430
rect 24278 70 24834 430
rect 24950 70 25506 430
rect 25622 70 26178 430
rect 26294 70 26850 430
rect 26966 70 27522 430
rect 27638 70 28194 430
rect 28310 70 28866 430
rect 28982 70 29538 430
rect 29654 70 30210 430
rect 30326 70 30882 430
rect 30998 70 31554 430
rect 31670 70 32226 430
rect 32342 70 32898 430
rect 33014 70 33570 430
rect 33686 70 34242 430
rect 34358 70 34914 430
rect 35030 70 35586 430
rect 35702 70 36258 430
rect 36374 70 36594 430
rect 36710 70 37266 430
rect 37382 70 37938 430
rect 38054 70 38610 430
rect 38726 70 39282 430
rect 39398 70 39954 430
rect 40070 70 40626 430
rect 40742 70 41298 430
rect 41414 70 41970 430
rect 42086 70 42642 430
rect 42758 70 43314 430
rect 43430 70 43986 430
rect 44102 70 44658 430
rect 44774 70 45330 430
rect 45446 70 46002 430
rect 46118 70 46674 430
rect 46790 70 47346 430
rect 47462 70 48018 430
rect 48134 70 48690 430
rect 48806 70 49362 430
rect 49478 70 50034 430
rect 50150 70 50706 430
rect 50822 70 51378 430
rect 51494 70 52050 430
rect 52166 70 52722 430
rect 52838 70 53394 430
rect 53510 70 54066 430
rect 54182 70 54402 430
rect 54518 70 55074 430
rect 55190 70 55746 430
rect 55862 70 56418 430
rect 56534 70 57090 430
rect 57206 70 57762 430
rect 57878 70 58434 430
rect 58550 70 59106 430
rect 59222 70 59778 430
rect 59894 70 60450 430
rect 60566 70 61122 430
rect 61238 70 61794 430
rect 61910 70 62466 430
rect 62582 70 63138 430
rect 63254 70 63810 430
rect 63926 70 64482 430
rect 64598 70 65154 430
rect 65270 70 65826 430
rect 65942 70 66498 430
rect 66614 70 67170 430
rect 67286 70 67842 430
rect 67958 70 68514 430
rect 68630 70 69186 430
rect 69302 70 69858 430
rect 69974 70 70530 430
rect 70646 70 71202 430
rect 71318 70 71874 430
rect 71990 70 72546 430
rect 72662 70 72882 430
rect 72998 70 73554 430
rect 73670 70 74226 430
rect 74342 70 74898 430
rect 75014 70 75570 430
rect 75686 70 76242 430
rect 76358 70 76914 430
rect 77030 70 77586 430
rect 77702 70 78258 430
rect 78374 70 78930 430
rect 79046 70 79602 430
rect 79718 70 80274 430
rect 80390 70 80946 430
rect 81062 70 81618 430
rect 81734 70 82290 430
rect 82406 70 82962 430
rect 83078 70 83634 430
rect 83750 70 84306 430
rect 84422 70 84978 430
rect 85094 70 85650 430
rect 85766 70 86322 430
rect 86438 70 86994 430
rect 87110 70 87666 430
rect 87782 70 88338 430
rect 88454 70 89010 430
rect 89126 70 89682 430
rect 89798 70 90354 430
rect 90470 70 90690 430
rect 90806 70 91362 430
rect 91478 70 92034 430
rect 92150 70 92706 430
rect 92822 70 93378 430
rect 93494 70 94050 430
rect 94166 70 94722 430
rect 94838 70 95394 430
rect 95510 70 96066 430
rect 96182 70 96738 430
rect 96854 70 97410 430
rect 97526 70 98082 430
rect 98198 70 98754 430
rect 98870 70 99162 430
rect 14 9 99162 70
<< metal3 >>
rect 99600 99792 99900 99848
rect 100 99456 400 99512
rect 99600 99120 99900 99176
rect 100 98784 400 98840
rect 99600 98448 99900 98504
rect 100 98112 400 98168
rect 99600 97776 99900 97832
rect 100 97440 400 97496
rect 99600 97104 99900 97160
rect 100 96768 400 96824
rect 99600 96432 99900 96488
rect 100 96096 400 96152
rect 99600 95760 99900 95816
rect 100 95424 400 95480
rect 99600 95088 99900 95144
rect 100 94752 400 94808
rect 99600 94416 99900 94472
rect 100 94080 400 94136
rect 99600 93744 99900 93800
rect 100 93408 400 93464
rect 99600 93072 99900 93128
rect 100 92736 400 92792
rect 99600 92400 99900 92456
rect 100 92064 400 92120
rect 99600 91728 99900 91784
rect 100 91392 400 91448
rect 99600 91056 99900 91112
rect 100 90720 400 90776
rect 100 90384 400 90440
rect 99600 90384 99900 90440
rect 100 89712 400 89768
rect 99600 89712 99900 89768
rect 100 89040 400 89096
rect 99600 89040 99900 89096
rect 100 88368 400 88424
rect 99600 88368 99900 88424
rect 100 87696 400 87752
rect 99600 87696 99900 87752
rect 100 87024 400 87080
rect 99600 87024 99900 87080
rect 100 86352 400 86408
rect 99600 86352 99900 86408
rect 100 85680 400 85736
rect 99600 85680 99900 85736
rect 100 85008 400 85064
rect 99600 85008 99900 85064
rect 100 84336 400 84392
rect 99600 84336 99900 84392
rect 100 83664 400 83720
rect 99600 83664 99900 83720
rect 100 82992 400 83048
rect 99600 82992 99900 83048
rect 100 82320 400 82376
rect 99600 82320 99900 82376
rect 100 81648 400 81704
rect 99600 81648 99900 81704
rect 99600 81312 99900 81368
rect 100 80976 400 81032
rect 99600 80640 99900 80696
rect 100 80304 400 80360
rect 99600 79968 99900 80024
rect 100 79632 400 79688
rect 99600 79296 99900 79352
rect 100 78960 400 79016
rect 99600 78624 99900 78680
rect 100 78288 400 78344
rect 99600 77952 99900 78008
rect 100 77616 400 77672
rect 99600 77280 99900 77336
rect 100 76944 400 77000
rect 99600 76608 99900 76664
rect 100 76272 400 76328
rect 99600 75936 99900 75992
rect 100 75600 400 75656
rect 99600 75264 99900 75320
rect 100 74928 400 74984
rect 99600 74592 99900 74648
rect 100 74256 400 74312
rect 99600 73920 99900 73976
rect 100 73584 400 73640
rect 99600 73248 99900 73304
rect 100 72912 400 72968
rect 100 72576 400 72632
rect 99600 72576 99900 72632
rect 100 71904 400 71960
rect 99600 71904 99900 71960
rect 100 71232 400 71288
rect 99600 71232 99900 71288
rect 100 70560 400 70616
rect 99600 70560 99900 70616
rect 100 69888 400 69944
rect 99600 69888 99900 69944
rect 100 69216 400 69272
rect 99600 69216 99900 69272
rect 100 68544 400 68600
rect 99600 68544 99900 68600
rect 100 67872 400 67928
rect 99600 67872 99900 67928
rect 100 67200 400 67256
rect 99600 67200 99900 67256
rect 100 66528 400 66584
rect 99600 66528 99900 66584
rect 100 65856 400 65912
rect 99600 65856 99900 65912
rect 100 65184 400 65240
rect 99600 65184 99900 65240
rect 100 64512 400 64568
rect 99600 64512 99900 64568
rect 100 63840 400 63896
rect 99600 63840 99900 63896
rect 99600 63504 99900 63560
rect 100 63168 400 63224
rect 99600 62832 99900 62888
rect 100 62496 400 62552
rect 99600 62160 99900 62216
rect 100 61824 400 61880
rect 99600 61488 99900 61544
rect 100 61152 400 61208
rect 99600 60816 99900 60872
rect 100 60480 400 60536
rect 99600 60144 99900 60200
rect 100 59808 400 59864
rect 99600 59472 99900 59528
rect 100 59136 400 59192
rect 99600 58800 99900 58856
rect 100 58464 400 58520
rect 99600 58128 99900 58184
rect 100 57792 400 57848
rect 99600 57456 99900 57512
rect 100 57120 400 57176
rect 99600 56784 99900 56840
rect 100 56448 400 56504
rect 99600 56112 99900 56168
rect 100 55776 400 55832
rect 99600 55440 99900 55496
rect 100 55104 400 55160
rect 99600 54768 99900 54824
rect 100 54432 400 54488
rect 100 54096 400 54152
rect 99600 54096 99900 54152
rect 100 53424 400 53480
rect 99600 53424 99900 53480
rect 100 52752 400 52808
rect 99600 52752 99900 52808
rect 100 52080 400 52136
rect 99600 52080 99900 52136
rect 100 51408 400 51464
rect 99600 51408 99900 51464
rect 100 50736 400 50792
rect 99600 50736 99900 50792
rect 100 50064 400 50120
rect 99600 50064 99900 50120
rect 100 49392 400 49448
rect 99600 49392 99900 49448
rect 100 48720 400 48776
rect 99600 48720 99900 48776
rect 100 48048 400 48104
rect 99600 48048 99900 48104
rect 100 47376 400 47432
rect 99600 47376 99900 47432
rect 100 46704 400 46760
rect 99600 46704 99900 46760
rect 100 46032 400 46088
rect 99600 46032 99900 46088
rect 100 45360 400 45416
rect 99600 45360 99900 45416
rect 99600 45024 99900 45080
rect 100 44688 400 44744
rect 99600 44352 99900 44408
rect 100 44016 400 44072
rect 99600 43680 99900 43736
rect 100 43344 400 43400
rect 99600 43008 99900 43064
rect 100 42672 400 42728
rect 99600 42336 99900 42392
rect 100 42000 400 42056
rect 99600 41664 99900 41720
rect 100 41328 400 41384
rect 99600 40992 99900 41048
rect 100 40656 400 40712
rect 99600 40320 99900 40376
rect 100 39984 400 40040
rect 99600 39648 99900 39704
rect 100 39312 400 39368
rect 99600 38976 99900 39032
rect 100 38640 400 38696
rect 99600 38304 99900 38360
rect 100 37968 400 38024
rect 99600 37632 99900 37688
rect 100 37296 400 37352
rect 99600 36960 99900 37016
rect 100 36624 400 36680
rect 100 36288 400 36344
rect 99600 36288 99900 36344
rect 100 35616 400 35672
rect 99600 35616 99900 35672
rect 100 34944 400 35000
rect 99600 34944 99900 35000
rect 100 34272 400 34328
rect 99600 34272 99900 34328
rect 100 33600 400 33656
rect 99600 33600 99900 33656
rect 100 32928 400 32984
rect 99600 32928 99900 32984
rect 100 32256 400 32312
rect 99600 32256 99900 32312
rect 100 31584 400 31640
rect 99600 31584 99900 31640
rect 100 30912 400 30968
rect 99600 30912 99900 30968
rect 100 30240 400 30296
rect 99600 30240 99900 30296
rect 100 29568 400 29624
rect 99600 29568 99900 29624
rect 100 28896 400 28952
rect 99600 28896 99900 28952
rect 100 28224 400 28280
rect 99600 28224 99900 28280
rect 100 27552 400 27608
rect 99600 27552 99900 27608
rect 99600 27216 99900 27272
rect 100 26880 400 26936
rect 99600 26544 99900 26600
rect 100 26208 400 26264
rect 99600 25872 99900 25928
rect 100 25536 400 25592
rect 99600 25200 99900 25256
rect 100 24864 400 24920
rect 99600 24528 99900 24584
rect 100 24192 400 24248
rect 99600 23856 99900 23912
rect 100 23520 400 23576
rect 99600 23184 99900 23240
rect 100 22848 400 22904
rect 99600 22512 99900 22568
rect 100 22176 400 22232
rect 99600 21840 99900 21896
rect 100 21504 400 21560
rect 99600 21168 99900 21224
rect 100 20832 400 20888
rect 99600 20496 99900 20552
rect 100 20160 400 20216
rect 99600 19824 99900 19880
rect 100 19488 400 19544
rect 99600 19152 99900 19208
rect 100 18816 400 18872
rect 99600 18480 99900 18536
rect 100 18144 400 18200
rect 100 17808 400 17864
rect 99600 17808 99900 17864
rect 100 17136 400 17192
rect 99600 17136 99900 17192
rect 100 16464 400 16520
rect 99600 16464 99900 16520
rect 100 15792 400 15848
rect 99600 15792 99900 15848
rect 100 15120 400 15176
rect 99600 15120 99900 15176
rect 100 14448 400 14504
rect 99600 14448 99900 14504
rect 100 13776 400 13832
rect 99600 13776 99900 13832
rect 100 13104 400 13160
rect 99600 13104 99900 13160
rect 100 12432 400 12488
rect 99600 12432 99900 12488
rect 100 11760 400 11816
rect 99600 11760 99900 11816
rect 100 11088 400 11144
rect 99600 11088 99900 11144
rect 100 10416 400 10472
rect 99600 10416 99900 10472
rect 100 9744 400 9800
rect 99600 9744 99900 9800
rect 100 9072 400 9128
rect 99600 9072 99900 9128
rect 99600 8736 99900 8792
rect 100 8400 400 8456
rect 99600 8064 99900 8120
rect 100 7728 400 7784
rect 99600 7392 99900 7448
rect 100 7056 400 7112
rect 99600 6720 99900 6776
rect 100 6384 400 6440
rect 99600 6048 99900 6104
rect 100 5712 400 5768
rect 99600 5376 99900 5432
rect 100 5040 400 5096
rect 99600 4704 99900 4760
rect 100 4368 400 4424
rect 99600 4032 99900 4088
rect 100 3696 400 3752
rect 99600 3360 99900 3416
rect 100 3024 400 3080
rect 99600 2688 99900 2744
rect 100 2352 400 2408
rect 99600 2016 99900 2072
rect 100 1680 400 1736
rect 99600 1344 99900 1400
rect 100 1008 400 1064
rect 99600 672 99900 728
rect 100 336 400 392
rect 99600 0 99900 56
<< obsm3 >>
rect 9 99090 99570 99162
rect 9 98870 99600 99090
rect 9 98754 70 98870
rect 430 98754 99600 98870
rect 9 98534 99600 98754
rect 9 98418 99570 98534
rect 9 98198 99600 98418
rect 9 98082 70 98198
rect 430 98082 99600 98198
rect 9 97862 99600 98082
rect 9 97746 99570 97862
rect 9 97526 99600 97746
rect 9 97410 70 97526
rect 430 97410 99600 97526
rect 9 97190 99600 97410
rect 9 97074 99570 97190
rect 9 96854 99600 97074
rect 9 96738 70 96854
rect 430 96738 99600 96854
rect 9 96518 99600 96738
rect 9 96402 99570 96518
rect 9 96182 99600 96402
rect 9 96066 70 96182
rect 430 96066 99600 96182
rect 9 95846 99600 96066
rect 9 95730 99570 95846
rect 9 95510 99600 95730
rect 9 95394 70 95510
rect 430 95394 99600 95510
rect 9 95174 99600 95394
rect 9 95058 99570 95174
rect 9 94838 99600 95058
rect 9 94722 70 94838
rect 430 94722 99600 94838
rect 9 94502 99600 94722
rect 9 94386 99570 94502
rect 9 94166 99600 94386
rect 9 94050 70 94166
rect 430 94050 99600 94166
rect 9 93830 99600 94050
rect 9 93714 99570 93830
rect 9 93494 99600 93714
rect 9 93378 70 93494
rect 430 93378 99600 93494
rect 9 93158 99600 93378
rect 9 93042 99570 93158
rect 9 92822 99600 93042
rect 9 92706 70 92822
rect 430 92706 99600 92822
rect 9 92486 99600 92706
rect 9 92370 99570 92486
rect 9 92150 99600 92370
rect 9 92034 70 92150
rect 430 92034 99600 92150
rect 9 91814 99600 92034
rect 9 91698 99570 91814
rect 9 91478 99600 91698
rect 9 91362 70 91478
rect 430 91362 99600 91478
rect 9 91142 99600 91362
rect 9 91026 99570 91142
rect 9 90806 99600 91026
rect 9 90690 70 90806
rect 430 90690 99600 90806
rect 9 90470 99600 90690
rect 9 90354 70 90470
rect 430 90354 99570 90470
rect 9 89798 99600 90354
rect 9 89682 70 89798
rect 430 89682 99570 89798
rect 9 89126 99600 89682
rect 9 89010 70 89126
rect 430 89010 99570 89126
rect 9 88454 99600 89010
rect 9 88338 70 88454
rect 430 88338 99570 88454
rect 9 87782 99600 88338
rect 9 87666 70 87782
rect 430 87666 99570 87782
rect 9 87110 99600 87666
rect 9 86994 70 87110
rect 430 86994 99570 87110
rect 9 86438 99600 86994
rect 9 86322 70 86438
rect 430 86322 99570 86438
rect 9 85766 99600 86322
rect 9 85650 70 85766
rect 430 85650 99570 85766
rect 9 85094 99600 85650
rect 9 84978 70 85094
rect 430 84978 99570 85094
rect 9 84422 99600 84978
rect 9 84306 70 84422
rect 430 84306 99570 84422
rect 9 83750 99600 84306
rect 9 83634 70 83750
rect 430 83634 99570 83750
rect 9 83078 99600 83634
rect 9 82962 70 83078
rect 430 82962 99570 83078
rect 9 82406 99600 82962
rect 9 82290 70 82406
rect 430 82290 99570 82406
rect 9 81734 99600 82290
rect 9 81618 70 81734
rect 430 81618 99570 81734
rect 9 81398 99600 81618
rect 9 81282 99570 81398
rect 9 81062 99600 81282
rect 9 80946 70 81062
rect 430 80946 99600 81062
rect 9 80726 99600 80946
rect 9 80610 99570 80726
rect 9 80390 99600 80610
rect 9 80274 70 80390
rect 430 80274 99600 80390
rect 9 80054 99600 80274
rect 9 79938 99570 80054
rect 9 79718 99600 79938
rect 9 79602 70 79718
rect 430 79602 99600 79718
rect 9 79382 99600 79602
rect 9 79266 99570 79382
rect 9 79046 99600 79266
rect 9 78930 70 79046
rect 430 78930 99600 79046
rect 9 78710 99600 78930
rect 9 78594 99570 78710
rect 9 78374 99600 78594
rect 9 78258 70 78374
rect 430 78258 99600 78374
rect 9 78038 99600 78258
rect 9 77922 99570 78038
rect 9 77702 99600 77922
rect 9 77586 70 77702
rect 430 77586 99600 77702
rect 9 77366 99600 77586
rect 9 77250 99570 77366
rect 9 77030 99600 77250
rect 9 76914 70 77030
rect 430 76914 99600 77030
rect 9 76694 99600 76914
rect 9 76578 99570 76694
rect 9 76358 99600 76578
rect 9 76242 70 76358
rect 430 76242 99600 76358
rect 9 76022 99600 76242
rect 9 75906 99570 76022
rect 9 75686 99600 75906
rect 9 75570 70 75686
rect 430 75570 99600 75686
rect 9 75350 99600 75570
rect 9 75234 99570 75350
rect 9 75014 99600 75234
rect 9 74898 70 75014
rect 430 74898 99600 75014
rect 9 74678 99600 74898
rect 9 74562 99570 74678
rect 9 74342 99600 74562
rect 9 74226 70 74342
rect 430 74226 99600 74342
rect 9 74006 99600 74226
rect 9 73890 99570 74006
rect 9 73670 99600 73890
rect 9 73554 70 73670
rect 430 73554 99600 73670
rect 9 73334 99600 73554
rect 9 73218 99570 73334
rect 9 72998 99600 73218
rect 9 72882 70 72998
rect 430 72882 99600 72998
rect 9 72662 99600 72882
rect 9 72546 70 72662
rect 430 72546 99570 72662
rect 9 71990 99600 72546
rect 9 71874 70 71990
rect 430 71874 99570 71990
rect 9 71318 99600 71874
rect 9 71202 70 71318
rect 430 71202 99570 71318
rect 9 70646 99600 71202
rect 9 70530 70 70646
rect 430 70530 99570 70646
rect 9 69974 99600 70530
rect 9 69858 70 69974
rect 430 69858 99570 69974
rect 9 69302 99600 69858
rect 9 69186 70 69302
rect 430 69186 99570 69302
rect 9 68630 99600 69186
rect 9 68514 70 68630
rect 430 68514 99570 68630
rect 9 67958 99600 68514
rect 9 67842 70 67958
rect 430 67842 99570 67958
rect 9 67286 99600 67842
rect 9 67170 70 67286
rect 430 67170 99570 67286
rect 9 66614 99600 67170
rect 9 66498 70 66614
rect 430 66498 99570 66614
rect 9 65942 99600 66498
rect 9 65826 70 65942
rect 430 65826 99570 65942
rect 9 65270 99600 65826
rect 9 65154 70 65270
rect 430 65154 99570 65270
rect 9 64598 99600 65154
rect 9 64482 70 64598
rect 430 64482 99570 64598
rect 9 63926 99600 64482
rect 9 63810 70 63926
rect 430 63810 99570 63926
rect 9 63590 99600 63810
rect 9 63474 99570 63590
rect 9 63254 99600 63474
rect 9 63138 70 63254
rect 430 63138 99600 63254
rect 9 62918 99600 63138
rect 9 62802 99570 62918
rect 9 62582 99600 62802
rect 9 62466 70 62582
rect 430 62466 99600 62582
rect 9 62246 99600 62466
rect 9 62130 99570 62246
rect 9 61910 99600 62130
rect 9 61794 70 61910
rect 430 61794 99600 61910
rect 9 61574 99600 61794
rect 9 61458 99570 61574
rect 9 61238 99600 61458
rect 9 61122 70 61238
rect 430 61122 99600 61238
rect 9 60902 99600 61122
rect 9 60786 99570 60902
rect 9 60566 99600 60786
rect 9 60450 70 60566
rect 430 60450 99600 60566
rect 9 60230 99600 60450
rect 9 60114 99570 60230
rect 9 59894 99600 60114
rect 9 59778 70 59894
rect 430 59778 99600 59894
rect 9 59558 99600 59778
rect 9 59442 99570 59558
rect 9 59222 99600 59442
rect 9 59106 70 59222
rect 430 59106 99600 59222
rect 9 58886 99600 59106
rect 9 58770 99570 58886
rect 9 58550 99600 58770
rect 9 58434 70 58550
rect 430 58434 99600 58550
rect 9 58214 99600 58434
rect 9 58098 99570 58214
rect 9 57878 99600 58098
rect 9 57762 70 57878
rect 430 57762 99600 57878
rect 9 57542 99600 57762
rect 9 57426 99570 57542
rect 9 57206 99600 57426
rect 9 57090 70 57206
rect 430 57090 99600 57206
rect 9 56870 99600 57090
rect 9 56754 99570 56870
rect 9 56534 99600 56754
rect 9 56418 70 56534
rect 430 56418 99600 56534
rect 9 56198 99600 56418
rect 9 56082 99570 56198
rect 9 55862 99600 56082
rect 9 55746 70 55862
rect 430 55746 99600 55862
rect 9 55526 99600 55746
rect 9 55410 99570 55526
rect 9 55190 99600 55410
rect 9 55074 70 55190
rect 430 55074 99600 55190
rect 9 54854 99600 55074
rect 9 54738 99570 54854
rect 9 54518 99600 54738
rect 9 54402 70 54518
rect 430 54402 99600 54518
rect 9 54182 99600 54402
rect 9 54066 70 54182
rect 430 54066 99570 54182
rect 9 53510 99600 54066
rect 9 53394 70 53510
rect 430 53394 99570 53510
rect 9 52838 99600 53394
rect 9 52722 70 52838
rect 430 52722 99570 52838
rect 9 52166 99600 52722
rect 9 52050 70 52166
rect 430 52050 99570 52166
rect 9 51494 99600 52050
rect 9 51378 70 51494
rect 430 51378 99570 51494
rect 9 50822 99600 51378
rect 9 50706 70 50822
rect 430 50706 99570 50822
rect 9 50150 99600 50706
rect 9 50034 70 50150
rect 430 50034 99570 50150
rect 9 49478 99600 50034
rect 9 49362 70 49478
rect 430 49362 99570 49478
rect 9 48806 99600 49362
rect 9 48690 70 48806
rect 430 48690 99570 48806
rect 9 48134 99600 48690
rect 9 48018 70 48134
rect 430 48018 99570 48134
rect 9 47462 99600 48018
rect 9 47346 70 47462
rect 430 47346 99570 47462
rect 9 46790 99600 47346
rect 9 46674 70 46790
rect 430 46674 99570 46790
rect 9 46118 99600 46674
rect 9 46002 70 46118
rect 430 46002 99570 46118
rect 9 45446 99600 46002
rect 9 45330 70 45446
rect 430 45330 99570 45446
rect 9 45110 99600 45330
rect 9 44994 99570 45110
rect 9 44774 99600 44994
rect 9 44658 70 44774
rect 430 44658 99600 44774
rect 9 44438 99600 44658
rect 9 44322 99570 44438
rect 9 44102 99600 44322
rect 9 43986 70 44102
rect 430 43986 99600 44102
rect 9 43766 99600 43986
rect 9 43650 99570 43766
rect 9 43430 99600 43650
rect 9 43314 70 43430
rect 430 43314 99600 43430
rect 9 43094 99600 43314
rect 9 42978 99570 43094
rect 9 42758 99600 42978
rect 9 42642 70 42758
rect 430 42642 99600 42758
rect 9 42422 99600 42642
rect 9 42306 99570 42422
rect 9 42086 99600 42306
rect 9 41970 70 42086
rect 430 41970 99600 42086
rect 9 41750 99600 41970
rect 9 41634 99570 41750
rect 9 41414 99600 41634
rect 9 41298 70 41414
rect 430 41298 99600 41414
rect 9 41078 99600 41298
rect 9 40962 99570 41078
rect 9 40742 99600 40962
rect 9 40626 70 40742
rect 430 40626 99600 40742
rect 9 40406 99600 40626
rect 9 40290 99570 40406
rect 9 40070 99600 40290
rect 9 39954 70 40070
rect 430 39954 99600 40070
rect 9 39734 99600 39954
rect 9 39618 99570 39734
rect 9 39398 99600 39618
rect 9 39282 70 39398
rect 430 39282 99600 39398
rect 9 39062 99600 39282
rect 9 38946 99570 39062
rect 9 38726 99600 38946
rect 9 38610 70 38726
rect 430 38610 99600 38726
rect 9 38390 99600 38610
rect 9 38274 99570 38390
rect 9 38054 99600 38274
rect 9 37938 70 38054
rect 430 37938 99600 38054
rect 9 37718 99600 37938
rect 9 37602 99570 37718
rect 9 37382 99600 37602
rect 9 37266 70 37382
rect 430 37266 99600 37382
rect 9 37046 99600 37266
rect 9 36930 99570 37046
rect 9 36710 99600 36930
rect 9 36594 70 36710
rect 430 36594 99600 36710
rect 9 36374 99600 36594
rect 9 36258 70 36374
rect 430 36258 99570 36374
rect 9 35702 99600 36258
rect 9 35586 70 35702
rect 430 35586 99570 35702
rect 9 35030 99600 35586
rect 9 34914 70 35030
rect 430 34914 99570 35030
rect 9 34358 99600 34914
rect 9 34242 70 34358
rect 430 34242 99570 34358
rect 9 33686 99600 34242
rect 9 33570 70 33686
rect 430 33570 99570 33686
rect 9 33014 99600 33570
rect 9 32898 70 33014
rect 430 32898 99570 33014
rect 9 32342 99600 32898
rect 9 32226 70 32342
rect 430 32226 99570 32342
rect 9 31670 99600 32226
rect 9 31554 70 31670
rect 430 31554 99570 31670
rect 9 30998 99600 31554
rect 9 30882 70 30998
rect 430 30882 99570 30998
rect 9 30326 99600 30882
rect 9 30210 70 30326
rect 430 30210 99570 30326
rect 9 29654 99600 30210
rect 9 29538 70 29654
rect 430 29538 99570 29654
rect 9 28982 99600 29538
rect 9 28866 70 28982
rect 430 28866 99570 28982
rect 9 28310 99600 28866
rect 9 28194 70 28310
rect 430 28194 99570 28310
rect 9 27638 99600 28194
rect 9 27522 70 27638
rect 430 27522 99570 27638
rect 9 27302 99600 27522
rect 9 27186 99570 27302
rect 9 26966 99600 27186
rect 9 26850 70 26966
rect 430 26850 99600 26966
rect 9 26630 99600 26850
rect 9 26514 99570 26630
rect 9 26294 99600 26514
rect 9 26178 70 26294
rect 430 26178 99600 26294
rect 9 25958 99600 26178
rect 9 25842 99570 25958
rect 9 25622 99600 25842
rect 9 25506 70 25622
rect 430 25506 99600 25622
rect 9 25286 99600 25506
rect 9 25170 99570 25286
rect 9 24950 99600 25170
rect 9 24834 70 24950
rect 430 24834 99600 24950
rect 9 24614 99600 24834
rect 9 24498 99570 24614
rect 9 24278 99600 24498
rect 9 24162 70 24278
rect 430 24162 99600 24278
rect 9 23942 99600 24162
rect 9 23826 99570 23942
rect 9 23606 99600 23826
rect 9 23490 70 23606
rect 430 23490 99600 23606
rect 9 23270 99600 23490
rect 9 23154 99570 23270
rect 9 22934 99600 23154
rect 9 22818 70 22934
rect 430 22818 99600 22934
rect 9 22598 99600 22818
rect 9 22482 99570 22598
rect 9 22262 99600 22482
rect 9 22146 70 22262
rect 430 22146 99600 22262
rect 9 21926 99600 22146
rect 9 21810 99570 21926
rect 9 21590 99600 21810
rect 9 21474 70 21590
rect 430 21474 99600 21590
rect 9 21254 99600 21474
rect 9 21138 99570 21254
rect 9 20918 99600 21138
rect 9 20802 70 20918
rect 430 20802 99600 20918
rect 9 20582 99600 20802
rect 9 20466 99570 20582
rect 9 20246 99600 20466
rect 9 20130 70 20246
rect 430 20130 99600 20246
rect 9 19910 99600 20130
rect 9 19794 99570 19910
rect 9 19574 99600 19794
rect 9 19458 70 19574
rect 430 19458 99600 19574
rect 9 19238 99600 19458
rect 9 19122 99570 19238
rect 9 18902 99600 19122
rect 9 18786 70 18902
rect 430 18786 99600 18902
rect 9 18566 99600 18786
rect 9 18450 99570 18566
rect 9 18230 99600 18450
rect 9 18114 70 18230
rect 430 18114 99600 18230
rect 9 17894 99600 18114
rect 9 17778 70 17894
rect 430 17778 99570 17894
rect 9 17222 99600 17778
rect 9 17106 70 17222
rect 430 17106 99570 17222
rect 9 16550 99600 17106
rect 9 16434 70 16550
rect 430 16434 99570 16550
rect 9 15878 99600 16434
rect 9 15762 70 15878
rect 430 15762 99570 15878
rect 9 15206 99600 15762
rect 9 15090 70 15206
rect 430 15090 99570 15206
rect 9 14534 99600 15090
rect 9 14418 70 14534
rect 430 14418 99570 14534
rect 9 13862 99600 14418
rect 9 13746 70 13862
rect 430 13746 99570 13862
rect 9 13190 99600 13746
rect 9 13074 70 13190
rect 430 13074 99570 13190
rect 9 12518 99600 13074
rect 9 12402 70 12518
rect 430 12402 99570 12518
rect 9 11846 99600 12402
rect 9 11730 70 11846
rect 430 11730 99570 11846
rect 9 11174 99600 11730
rect 9 11058 70 11174
rect 430 11058 99570 11174
rect 9 10502 99600 11058
rect 9 10386 70 10502
rect 430 10386 99570 10502
rect 9 9830 99600 10386
rect 9 9714 70 9830
rect 430 9714 99570 9830
rect 9 9158 99600 9714
rect 9 9042 70 9158
rect 430 9042 99570 9158
rect 9 8822 99600 9042
rect 9 8706 99570 8822
rect 9 8486 99600 8706
rect 9 8370 70 8486
rect 430 8370 99600 8486
rect 9 8150 99600 8370
rect 9 8034 99570 8150
rect 9 7814 99600 8034
rect 9 7698 70 7814
rect 430 7698 99600 7814
rect 9 7478 99600 7698
rect 9 7362 99570 7478
rect 9 7142 99600 7362
rect 9 7026 70 7142
rect 430 7026 99600 7142
rect 9 6806 99600 7026
rect 9 6690 99570 6806
rect 9 6470 99600 6690
rect 9 6354 70 6470
rect 430 6354 99600 6470
rect 9 6134 99600 6354
rect 9 6018 99570 6134
rect 9 5798 99600 6018
rect 9 5682 70 5798
rect 430 5682 99600 5798
rect 9 5462 99600 5682
rect 9 5346 99570 5462
rect 9 5126 99600 5346
rect 9 5010 70 5126
rect 430 5010 99600 5126
rect 9 4790 99600 5010
rect 9 4674 99570 4790
rect 9 4454 99600 4674
rect 9 4338 70 4454
rect 430 4338 99600 4454
rect 9 4118 99600 4338
rect 9 4002 99570 4118
rect 9 3782 99600 4002
rect 9 3666 70 3782
rect 430 3666 99600 3782
rect 9 3446 99600 3666
rect 9 3330 99570 3446
rect 9 3110 99600 3330
rect 9 2994 70 3110
rect 430 2994 99600 3110
rect 9 2774 99600 2994
rect 9 2658 99570 2774
rect 9 2438 99600 2658
rect 9 2322 70 2438
rect 430 2322 99600 2438
rect 9 2102 99600 2322
rect 9 1986 99570 2102
rect 9 1766 99600 1986
rect 9 1650 70 1766
rect 430 1650 99600 1766
rect 9 1430 99600 1650
rect 9 1314 99570 1430
rect 9 1094 99600 1314
rect 9 978 70 1094
rect 430 978 99600 1094
rect 9 758 99600 978
rect 9 642 99570 758
rect 9 422 99600 642
rect 9 306 70 422
rect 430 306 99600 422
rect 9 86 99600 306
rect 9 14 99570 86
<< metal4 >>
rect 2224 1538 2384 98422
rect 9904 1538 10064 98422
rect 17584 1538 17744 98422
rect 25264 1538 25424 98422
rect 32944 1538 33104 98422
rect 40624 1538 40784 98422
rect 48304 1538 48464 98422
rect 55984 1538 56144 98422
rect 63664 1538 63824 98422
rect 71344 1538 71504 98422
rect 79024 1538 79184 98422
rect 86704 1538 86864 98422
rect 94384 1538 94544 98422
<< labels >>
rlabel metal2 s 98112 100 98168 400 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 5712 100 5768 400 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 99600 45024 99900 45080 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 100 21504 400 21560 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 32256 99600 32312 99900 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 99600 65856 99900 65912 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 27216 99600 27272 99900 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 100 10416 400 10472 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 99600 95760 99900 95816 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 100 33600 400 33656 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 35616 99600 35672 99900 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 9072 100 9128 400 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 23856 99600 23912 99900 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 28896 99600 28952 99900 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 100 9072 400 9128 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 100 24864 400 24920 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 99600 74592 99900 74648 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 2016 99600 2072 99900 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 62160 99600 62216 99900 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 25872 99600 25928 99900 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 100 3696 400 3752 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 44352 99600 44408 99900 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 100 81648 400 81704 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 42672 100 42728 400 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 100 28896 400 28952 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 67200 99600 67256 99900 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 57456 99600 57512 99900 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 30240 100 30296 400 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 99600 66528 99900 66584 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 100 34272 400 34328 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 92736 100 92792 400 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 100 34944 400 35000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 94416 99600 94472 99900 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 99600 13104 99900 13160 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 99600 59472 99900 59528 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 100 55104 400 55160 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 46704 99600 46760 99900 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 100 64512 400 64568 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 99600 36288 99900 36344 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 99600 34272 99900 34328 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 58800 99600 58856 99900 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 33600 99600 33656 99900 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 74256 100 74312 400 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 15792 99600 15848 99900 6 io_oeb[14]
port 44 nsew signal output
rlabel metal3 s 99600 36960 99900 37016 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 68544 100 68600 400 6 io_oeb[16]
port 46 nsew signal output
rlabel metal3 s 100 98784 400 98840 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 672 99600 728 99900 6 io_oeb[18]
port 48 nsew signal output
rlabel metal3 s 100 30240 400 30296 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 67872 100 67928 400 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 16464 99600 16520 99900 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 67872 99600 67928 99900 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 100 17808 400 17864 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 99600 41664 99900 41720 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 99600 99120 99900 99176 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 100 77616 400 77672 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 9744 99600 9800 99900 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 100 1008 400 1064 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 60144 99600 60200 99900 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 99600 73920 99900 73976 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 99600 86352 99900 86408 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 62496 100 62552 400 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 100 87696 400 87752 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 11088 99600 11144 99900 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 2688 99600 2744 99900 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 17136 99600 17192 99900 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 100 54096 400 54152 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 44688 100 44744 400 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 100 72912 400 72968 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 75936 99600 75992 99900 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 50736 100 50792 400 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 100 26880 400 26936 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 71232 99600 71288 99900 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 96432 99600 96488 99900 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 100 70560 400 70616 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 8736 99600 8792 99900 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 100 97440 400 97496 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 93744 99600 93800 99900 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 100 45360 400 45416 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 99600 93072 99900 93128 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 100 32256 400 32312 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 13104 100 13160 400 6 io_out[14]
port 82 nsew signal output
rlabel metal3 s 99600 77952 99900 78008 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 99600 23856 99900 23912 6 io_out[16]
port 84 nsew signal output
rlabel metal3 s 99600 65184 99900 65240 6 io_out[17]
port 85 nsew signal output
rlabel metal3 s 99600 89712 99900 89768 6 io_out[18]
port 86 nsew signal output
rlabel metal3 s 99600 78624 99900 78680 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 11760 100 11816 400 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 76944 100 77000 400 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 100 96096 400 96152 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 95424 100 95480 400 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 55776 100 55832 400 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 99600 11760 99900 11816 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 100 67872 400 67928 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 18480 99600 18536 99900 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 99600 672 99900 728 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 99600 56112 99900 56168 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 23520 100 23576 400 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 95760 99600 95816 99900 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 31584 100 31640 400 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 99600 88368 99900 88424 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 90720 100 90776 400 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 99600 75936 99900 75992 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 99120 99600 99176 99900 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 99600 67872 99900 67928 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 17808 99600 17864 99900 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 90384 100 90440 400 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 100 48720 400 48776 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 99600 10416 99900 10472 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 99600 62832 99900 62888 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 49392 99600 49448 99900 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 100 22848 400 22904 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 39648 99600 39704 99900 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 100 96768 400 96824 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 32256 100 32312 400 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 99600 40992 99900 41048 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 78624 99600 78680 99900 6 irq[2]
port 117 nsew signal output
rlabel metal3 s 99600 51408 99900 51464 6 la_data_in[0]
port 118 nsew signal input
rlabel metal3 s 99600 28896 99900 28952 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 43008 99600 43064 99900 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 14448 99600 14504 99900 6 la_data_in[102]
port 121 nsew signal input
rlabel metal3 s 99600 91728 99900 91784 6 la_data_in[103]
port 122 nsew signal input
rlabel metal3 s 100 74928 400 74984 6 la_data_in[104]
port 123 nsew signal input
rlabel metal3 s 99600 63504 99900 63560 6 la_data_in[105]
port 124 nsew signal input
rlabel metal3 s 99600 11088 99900 11144 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 53424 99600 53480 99900 6 la_data_in[107]
port 126 nsew signal input
rlabel metal3 s 99600 27216 99900 27272 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 70560 99600 70616 99900 6 la_data_in[109]
port 128 nsew signal input
rlabel metal3 s 100 76944 400 77000 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 3024 100 3080 400 6 la_data_in[110]
port 130 nsew signal input
rlabel metal3 s 99600 63840 99900 63896 6 la_data_in[111]
port 131 nsew signal input
rlabel metal3 s 100 78288 400 78344 6 la_data_in[112]
port 132 nsew signal input
rlabel metal3 s 99600 16464 99900 16520 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 73248 99600 73304 99900 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 24192 100 24248 400 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 44016 100 44072 400 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 38976 99600 39032 99900 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 79968 99600 80024 99900 6 la_data_in[118]
port 138 nsew signal input
rlabel metal3 s 99600 60816 99900 60872 6 la_data_in[119]
port 139 nsew signal input
rlabel metal3 s 100 71904 400 71960 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 66528 99600 66584 99900 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 97440 100 97496 400 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 3360 99600 3416 99900 6 la_data_in[122]
port 143 nsew signal input
rlabel metal3 s 99600 2016 99900 2072 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 7392 99600 7448 99900 6 la_data_in[124]
port 145 nsew signal input
rlabel metal3 s 100 25536 400 25592 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 76272 100 76328 400 6 la_data_in[126]
port 147 nsew signal input
rlabel metal3 s 100 53424 400 53480 6 la_data_in[127]
port 148 nsew signal input
rlabel metal3 s 100 44688 400 44744 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 89040 100 89096 400 6 la_data_in[13]
port 150 nsew signal input
rlabel metal3 s 99600 72576 99900 72632 6 la_data_in[14]
port 151 nsew signal input
rlabel metal3 s 100 15792 400 15848 6 la_data_in[15]
port 152 nsew signal input
rlabel metal3 s 99600 43008 99900 43064 6 la_data_in[16]
port 153 nsew signal input
rlabel metal3 s 100 40656 400 40712 6 la_data_in[17]
port 154 nsew signal input
rlabel metal3 s 99600 84336 99900 84392 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 75264 99600 75320 99900 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 24864 100 24920 400 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 0 99600 56 99900 6 la_data_in[20]
port 158 nsew signal input
rlabel metal3 s 100 3024 400 3080 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 66528 100 66584 400 6 la_data_in[22]
port 160 nsew signal input
rlabel metal3 s 99600 53424 99900 53480 6 la_data_in[23]
port 161 nsew signal input
rlabel metal3 s 99600 20496 99900 20552 6 la_data_in[24]
port 162 nsew signal input
rlabel metal3 s 100 65856 400 65912 6 la_data_in[25]
port 163 nsew signal input
rlabel metal3 s 99600 80640 99900 80696 6 la_data_in[26]
port 164 nsew signal input
rlabel metal3 s 100 7056 400 7112 6 la_data_in[27]
port 165 nsew signal input
rlabel metal3 s 99600 60144 99900 60200 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 71904 100 71960 400 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 79632 100 79688 400 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 94080 100 94136 400 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 34944 99600 35000 99900 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 72912 100 72968 400 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 41328 100 41384 400 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 45024 99600 45080 99900 6 la_data_in[34]
port 173 nsew signal input
rlabel metal3 s 100 82992 400 83048 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 77952 99600 78008 99900 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 97104 99600 97160 99900 6 la_data_in[37]
port 176 nsew signal input
rlabel metal3 s 99600 44352 99900 44408 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 1680 100 1736 400 6 la_data_in[39]
port 178 nsew signal input
rlabel metal3 s 100 51408 400 51464 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 20160 100 20216 400 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 26208 100 26264 400 6 la_data_in[41]
port 181 nsew signal input
rlabel metal3 s 99600 46032 99900 46088 6 la_data_in[42]
port 182 nsew signal input
rlabel metal3 s 99600 77280 99900 77336 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 31584 99600 31640 99900 6 la_data_in[44]
port 184 nsew signal input
rlabel metal3 s 100 17136 400 17192 6 la_data_in[45]
port 185 nsew signal input
rlabel metal3 s 100 54432 400 54488 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 67200 100 67256 400 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 69888 99600 69944 99900 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 19488 100 19544 400 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 34944 100 35000 400 6 la_data_in[4]
port 190 nsew signal input
rlabel metal3 s 100 1680 400 1736 6 la_data_in[50]
port 191 nsew signal input
rlabel metal3 s 100 99456 400 99512 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 95088 99600 95144 99900 6 la_data_in[52]
port 193 nsew signal input
rlabel metal3 s 99600 19824 99900 19880 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 12432 100 12488 400 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 47376 100 47432 400 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 336 100 392 400 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 74928 100 74984 400 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 82320 99600 82376 99900 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 87696 100 87752 400 6 la_data_in[59]
port 200 nsew signal input
rlabel metal3 s 100 42000 400 42056 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 6048 99600 6104 99900 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 20832 100 20888 400 6 la_data_in[61]
port 203 nsew signal input
rlabel metal3 s 99600 25200 99900 25256 6 la_data_in[62]
port 204 nsew signal input
rlabel metal3 s 100 55776 400 55832 6 la_data_in[63]
port 205 nsew signal input
rlabel metal3 s 99600 94416 99900 94472 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 87024 100 87080 400 6 la_data_in[65]
port 207 nsew signal input
rlabel metal3 s 100 93408 400 93464 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 40320 99600 40376 99900 6 la_data_in[67]
port 209 nsew signal input
rlabel metal3 s 100 24192 400 24248 6 la_data_in[68]
port 210 nsew signal input
rlabel metal3 s 99600 73248 99900 73304 6 la_data_in[69]
port 211 nsew signal input
rlabel metal3 s 99600 40320 99900 40376 6 la_data_in[6]
port 212 nsew signal input
rlabel metal3 s 99600 25872 99900 25928 6 la_data_in[70]
port 213 nsew signal input
rlabel metal3 s 99600 19152 99900 19208 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 23184 99600 23240 99900 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 99456 100 99512 400 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 49392 100 49448 400 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 39312 100 39368 400 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 48720 100 48776 400 6 la_data_in[76]
port 219 nsew signal input
rlabel metal3 s 99600 64512 99900 64568 6 la_data_in[77]
port 220 nsew signal input
rlabel metal3 s 99600 79968 99900 80024 6 la_data_in[78]
port 221 nsew signal input
rlabel metal3 s 99600 28224 99900 28280 6 la_data_in[79]
port 222 nsew signal input
rlabel metal3 s 99600 31584 99900 31640 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 82320 100 82376 400 6 la_data_in[80]
port 224 nsew signal input
rlabel metal3 s 99600 32256 99900 32312 6 la_data_in[81]
port 225 nsew signal input
rlabel metal3 s 100 44016 400 44072 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 82992 99600 83048 99900 6 la_data_in[83]
port 227 nsew signal input
rlabel metal3 s 100 336 400 392 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 38304 99600 38360 99900 6 la_data_in[85]
port 229 nsew signal input
rlabel metal3 s 99600 71232 99900 71288 6 la_data_in[86]
port 230 nsew signal input
rlabel metal3 s 100 50064 400 50120 6 la_data_in[87]
port 231 nsew signal input
rlabel metal3 s 100 60480 400 60536 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 32928 99600 32984 99900 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 21840 99600 21896 99900 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 56784 99600 56840 99900 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 1344 99600 1400 99900 6 la_data_in[91]
port 236 nsew signal input
rlabel metal3 s 99600 2688 99900 2744 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 35616 100 35672 400 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 39984 100 40040 400 6 la_data_in[94]
port 239 nsew signal input
rlabel metal3 s 99600 9072 99900 9128 6 la_data_in[95]
port 240 nsew signal input
rlabel metal3 s 100 35616 400 35672 6 la_data_in[96]
port 241 nsew signal input
rlabel metal3 s 100 87024 400 87080 6 la_data_in[97]
port 242 nsew signal input
rlabel metal3 s 99600 47376 99900 47432 6 la_data_in[98]
port 243 nsew signal input
rlabel metal3 s 100 67200 400 67256 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 17808 100 17864 400 6 la_data_in[9]
port 245 nsew signal input
rlabel metal3 s 100 62496 400 62552 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 92400 99600 92456 99900 6 la_data_out[100]
port 247 nsew signal output
rlabel metal3 s 100 86352 400 86408 6 la_data_out[101]
port 248 nsew signal output
rlabel metal3 s 100 8400 400 8456 6 la_data_out[102]
port 249 nsew signal output
rlabel metal3 s 99600 37632 99900 37688 6 la_data_out[103]
port 250 nsew signal output
rlabel metal3 s 99600 54768 99900 54824 6 la_data_out[104]
port 251 nsew signal output
rlabel metal3 s 100 31584 400 31640 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 21168 99600 21224 99900 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 65856 100 65912 400 6 la_data_out[107]
port 254 nsew signal output
rlabel metal3 s 100 78960 400 79016 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 50736 99600 50792 99900 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 59472 99600 59528 99900 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 15792 100 15848 400 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 72576 99600 72632 99900 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 90384 99600 90440 99900 6 la_data_out[112]
port 260 nsew signal output
rlabel metal3 s 100 7728 400 7784 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 40992 99600 41048 99900 6 la_data_out[114]
port 262 nsew signal output
rlabel metal3 s 99600 87696 99900 87752 6 la_data_out[115]
port 263 nsew signal output
rlabel metal3 s 99600 23184 99900 23240 6 la_data_out[116]
port 264 nsew signal output
rlabel metal3 s 100 23520 400 23576 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 37968 100 38024 400 6 la_data_out[118]
port 266 nsew signal output
rlabel metal3 s 100 36288 400 36344 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 57120 100 57176 400 6 la_data_out[11]
port 268 nsew signal output
rlabel metal3 s 99600 4032 99900 4088 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 15120 99600 15176 99900 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 91728 99600 91784 99900 6 la_data_out[122]
port 271 nsew signal output
rlabel metal3 s 100 79632 400 79688 6 la_data_out[123]
port 272 nsew signal output
rlabel metal3 s 100 32928 400 32984 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 91392 100 91448 400 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 57792 100 57848 400 6 la_data_out[126]
port 275 nsew signal output
rlabel metal3 s 100 59808 400 59864 6 la_data_out[127]
port 276 nsew signal output
rlabel metal3 s 99600 89040 99900 89096 6 la_data_out[12]
port 277 nsew signal output
rlabel metal3 s 99600 45360 99900 45416 6 la_data_out[13]
port 278 nsew signal output
rlabel metal3 s 100 38640 400 38696 6 la_data_out[14]
port 279 nsew signal output
rlabel metal3 s 99600 50064 99900 50120 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 98784 100 98840 400 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 6720 99600 6776 99900 6 la_data_out[17]
port 282 nsew signal output
rlabel metal3 s 99600 17808 99900 17864 6 la_data_out[18]
port 283 nsew signal output
rlabel metal3 s 100 63840 400 63896 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 5376 99600 5432 99900 6 la_data_out[1]
port 285 nsew signal output
rlabel metal3 s 99600 97104 99900 97160 6 la_data_out[20]
port 286 nsew signal output
rlabel metal3 s 100 20160 400 20216 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 64512 99600 64568 99900 6 la_data_out[22]
port 288 nsew signal output
rlabel metal3 s 99600 38304 99900 38360 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 46032 100 46088 400 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 54768 99600 54824 99900 6 la_data_out[25]
port 291 nsew signal output
rlabel metal3 s 100 19488 400 19544 6 la_data_out[26]
port 292 nsew signal output
rlabel metal3 s 99600 46704 99900 46760 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 15120 100 15176 400 6 la_data_out[28]
port 294 nsew signal output
rlabel metal3 s 100 92064 400 92120 6 la_data_out[29]
port 295 nsew signal output
rlabel metal3 s 99600 15120 99900 15176 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 46704 100 46760 400 6 la_data_out[30]
port 297 nsew signal output
rlabel metal3 s 100 29568 400 29624 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 19824 99600 19880 99900 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 56112 99600 56168 99900 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 96768 100 96824 400 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 87696 99600 87752 99900 6 la_data_out[35]
port 302 nsew signal output
rlabel metal3 s 100 74256 400 74312 6 la_data_out[36]
port 303 nsew signal output
rlabel metal3 s 100 47376 400 47432 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 79296 99600 79352 99900 6 la_data_out[38]
port 305 nsew signal output
rlabel metal3 s 99600 27552 99900 27608 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 36960 99600 37016 99900 6 la_data_out[3]
port 307 nsew signal output
rlabel metal3 s 100 63168 400 63224 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 56448 100 56504 400 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 29568 99600 29624 99900 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 26544 99600 26600 99900 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 84336 100 84392 400 6 la_data_out[44]
port 312 nsew signal output
rlabel metal3 s 99600 3360 99900 3416 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 98448 99600 98504 99900 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 34272 99600 34328 99900 6 la_data_out[47]
port 315 nsew signal output
rlabel metal3 s 100 11760 400 11816 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 7056 100 7112 400 6 la_data_out[49]
port 317 nsew signal output
rlabel metal3 s 100 46704 400 46760 6 la_data_out[4]
port 318 nsew signal output
rlabel metal3 s 100 56448 400 56504 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 30912 100 30968 400 6 la_data_out[51]
port 320 nsew signal output
rlabel metal3 s 100 75600 400 75656 6 la_data_out[52]
port 321 nsew signal output
rlabel metal3 s 99600 50736 99900 50792 6 la_data_out[53]
port 322 nsew signal output
rlabel metal3 s 100 61152 400 61208 6 la_data_out[54]
port 323 nsew signal output
rlabel metal3 s 99600 48048 99900 48104 6 la_data_out[55]
port 324 nsew signal output
rlabel metal3 s 100 5040 400 5096 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 52752 100 52808 400 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 93072 99600 93128 99900 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 76608 99600 76664 99900 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 47376 99600 47432 99900 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 13776 100 13832 400 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 78960 100 79016 400 6 la_data_out[61]
port 331 nsew signal output
rlabel metal3 s 100 85008 400 85064 6 la_data_out[62]
port 332 nsew signal output
rlabel metal3 s 99600 54096 99900 54152 6 la_data_out[63]
port 333 nsew signal output
rlabel metal3 s 99600 22512 99900 22568 6 la_data_out[64]
port 334 nsew signal output
rlabel metal3 s 99600 13776 99900 13832 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 48048 100 48104 400 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 71232 100 71288 400 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 36624 100 36680 400 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 89712 99600 89768 99900 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 54432 100 54488 400 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 37632 99600 37688 99900 6 la_data_out[70]
port 341 nsew signal output
rlabel metal3 s 100 94080 400 94136 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 26880 100 26936 400 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 48720 99600 48776 99900 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 50064 100 50120 400 6 la_data_out[74]
port 345 nsew signal output
rlabel metal3 s 99600 9744 99900 9800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 94752 100 94808 400 6 la_data_out[76]
port 347 nsew signal output
rlabel metal3 s 99600 21840 99900 21896 6 la_data_out[77]
port 348 nsew signal output
rlabel metal3 s 99600 17136 99900 17192 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 37296 100 37352 400 6 la_data_out[79]
port 350 nsew signal output
rlabel metal3 s 100 91392 400 91448 6 la_data_out[7]
port 351 nsew signal output
rlabel metal3 s 100 12432 400 12488 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 20496 99600 20552 99900 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 81648 100 81704 400 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 13104 99600 13160 99900 6 la_data_out[83]
port 355 nsew signal output
rlabel metal3 s 100 18144 400 18200 6 la_data_out[84]
port 356 nsew signal output
rlabel metal3 s 99600 0 99900 56 6 la_data_out[85]
port 357 nsew signal output
rlabel metal3 s 99600 52080 99900 52136 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 54096 99600 54152 99900 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 63840 100 63896 400 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 51408 99600 51464 99900 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 52080 99600 52136 99900 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 75600 100 75656 400 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 85008 100 85064 400 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 84336 99600 84392 99900 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 30912 99600 30968 99900 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 41664 99600 41720 99900 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 78288 100 78344 400 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 8064 99600 8120 99900 6 la_data_out[96]
port 369 nsew signal output
rlabel metal3 s 100 37296 400 37352 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 81648 99600 81704 99900 6 la_data_out[98]
port 371 nsew signal output
rlabel metal3 s 99600 1344 99900 1400 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 45360 100 45416 400 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 53424 100 53480 400 6 la_oenb[0]
port 374 nsew signal input
rlabel metal3 s 99600 98448 99900 98504 6 la_oenb[100]
port 375 nsew signal input
rlabel metal3 s 100 83664 400 83720 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 83664 99600 83720 99900 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 25536 100 25592 400 6 la_oenb[103]
port 378 nsew signal input
rlabel metal3 s 99600 58128 99900 58184 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 45360 99600 45416 99900 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 97776 99600 97832 99900 6 la_oenb[106]
port 381 nsew signal input
rlabel metal3 s 99600 56784 99900 56840 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 65184 99600 65240 99900 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 77280 99600 77336 99900 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 40656 100 40712 400 6 la_oenb[10]
port 385 nsew signal input
rlabel metal3 s 99600 76608 99900 76664 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 73584 100 73640 400 6 la_oenb[111]
port 387 nsew signal input
rlabel metal3 s 100 52080 400 52136 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 18816 100 18872 400 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 58128 99600 58184 99900 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 58464 100 58520 400 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 52080 100 52136 400 6 la_oenb[116]
port 392 nsew signal input
rlabel metal3 s 99600 95088 99900 95144 6 la_oenb[117]
port 393 nsew signal input
rlabel metal3 s 99600 39648 99900 39704 6 la_oenb[118]
port 394 nsew signal input
rlabel metal3 s 100 48048 400 48104 6 la_oenb[119]
port 395 nsew signal input
rlabel metal3 s 99600 57456 99900 57512 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 64512 100 64568 400 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 36288 100 36344 400 6 la_oenb[121]
port 398 nsew signal input
rlabel metal3 s 100 72576 400 72632 6 la_oenb[122]
port 399 nsew signal input
rlabel metal3 s 99600 82992 99900 83048 6 la_oenb[123]
port 400 nsew signal input
rlabel metal3 s 100 57792 400 57848 6 la_oenb[124]
port 401 nsew signal input
rlabel metal3 s 100 68544 400 68600 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 82992 100 83048 400 6 la_oenb[126]
port 403 nsew signal input
rlabel metal3 s 99600 26544 99900 26600 6 la_oenb[127]
port 404 nsew signal input
rlabel metal3 s 99600 69216 99900 69272 6 la_oenb[12]
port 405 nsew signal input
rlabel metal3 s 100 16464 400 16520 6 la_oenb[13]
port 406 nsew signal input
rlabel metal3 s 100 13776 400 13832 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 54096 100 54152 400 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 28896 100 28952 400 6 la_oenb[16]
port 409 nsew signal input
rlabel metal3 s 99600 18480 99900 18536 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 6384 100 6440 400 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 29568 100 29624 400 6 la_oenb[19]
port 412 nsew signal input
rlabel metal3 s 99600 15792 99900 15848 6 la_oenb[1]
port 413 nsew signal input
rlabel metal3 s 99600 93744 99900 93800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal3 s 99600 42336 99900 42392 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 10416 100 10472 400 6 la_oenb[22]
port 416 nsew signal input
rlabel metal3 s 100 30912 400 30968 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 70560 100 70616 400 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 87024 99600 87080 99900 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 65184 100 65240 400 6 la_oenb[26]
port 420 nsew signal input
rlabel metal3 s 99600 55440 99900 55496 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 99792 99600 99848 99900 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 88368 99600 88424 99900 6 la_oenb[29]
port 423 nsew signal input
rlabel metal3 s 100 4368 400 4424 6 la_oenb[2]
port 424 nsew signal input
rlabel metal3 s 100 46032 400 46088 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 27552 99600 27608 99900 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 33600 100 33656 400 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 10416 99600 10472 99900 6 la_oenb[33]
port 428 nsew signal input
rlabel metal3 s 99600 32928 99900 32984 6 la_oenb[34]
port 429 nsew signal input
rlabel metal3 s 99600 58800 99900 58856 6 la_oenb[35]
port 430 nsew signal input
rlabel metal3 s 100 13104 400 13160 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 77616 100 77672 400 6 la_oenb[37]
port 432 nsew signal input
rlabel metal3 s 99600 81648 99900 81704 6 la_oenb[38]
port 433 nsew signal input
rlabel metal3 s 100 66528 400 66584 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 91056 99600 91112 99900 6 la_oenb[3]
port 435 nsew signal input
rlabel metal3 s 100 85680 400 85736 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 93408 100 93464 400 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 4032 99600 4088 99900 6 la_oenb[42]
port 438 nsew signal input
rlabel metal3 s 100 84336 400 84392 6 la_oenb[43]
port 439 nsew signal input
rlabel metal3 s 99600 7392 99900 7448 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 18144 100 18200 400 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 27552 100 27608 400 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 96096 100 96152 400 6 la_oenb[47]
port 443 nsew signal input
rlabel metal3 s 99600 30912 99900 30968 6 la_oenb[48]
port 444 nsew signal input
rlabel metal3 s 99600 82320 99900 82376 6 la_oenb[49]
port 445 nsew signal input
rlabel metal3 s 100 69216 400 69272 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 46032 99600 46088 99900 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 30240 99600 30296 99900 6 la_oenb[51]
port 448 nsew signal input
rlabel metal3 s 100 49392 400 49448 6 la_oenb[52]
port 449 nsew signal input
rlabel metal3 s 99600 92400 99900 92456 6 la_oenb[53]
port 450 nsew signal input
rlabel metal3 s 100 73584 400 73640 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 24528 99600 24584 99900 6 la_oenb[55]
port 452 nsew signal input
rlabel metal3 s 100 14448 400 14504 6 la_oenb[56]
port 453 nsew signal input
rlabel metal3 s 99600 81312 99900 81368 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 69216 99600 69272 99900 6 la_oenb[58]
port 455 nsew signal input
rlabel metal3 s 100 92736 400 92792 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 80640 99600 80696 99900 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 85680 99600 85736 99900 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 86352 99600 86408 99900 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 59808 100 59864 400 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 52752 99600 52808 99900 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 3696 100 3752 400 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 1008 100 1064 400 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 89712 100 89768 400 6 la_oenb[66]
port 464 nsew signal input
rlabel metal3 s 100 41328 400 41384 6 la_oenb[67]
port 465 nsew signal input
rlabel metal3 s 99600 21168 99900 21224 6 la_oenb[68]
port 466 nsew signal input
rlabel metal3 s 100 52752 400 52808 6 la_oenb[69]
port 467 nsew signal input
rlabel metal3 s 100 69888 400 69944 6 la_oenb[6]
port 468 nsew signal input
rlabel metal3 s 100 95424 400 95480 6 la_oenb[70]
port 469 nsew signal input
rlabel metal3 s 100 43344 400 43400 6 la_oenb[71]
port 470 nsew signal input
rlabel metal3 s 100 36624 400 36680 6 la_oenb[72]
port 471 nsew signal input
rlabel metal3 s 100 28224 400 28280 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 50064 99600 50120 99900 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 92064 100 92120 400 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 43344 100 43400 400 6 la_oenb[76]
port 475 nsew signal input
rlabel metal3 s 100 80976 400 81032 6 la_oenb[77]
port 476 nsew signal input
rlabel metal3 s 99600 69888 99900 69944 6 la_oenb[78]
port 477 nsew signal input
rlabel metal3 s 99600 91056 99900 91112 6 la_oenb[79]
port 478 nsew signal input
rlabel metal3 s 100 58464 400 58520 6 la_oenb[7]
port 479 nsew signal input
rlabel metal3 s 100 71232 400 71288 6 la_oenb[80]
port 480 nsew signal input
rlabel metal3 s 99600 12432 99900 12488 6 la_oenb[81]
port 481 nsew signal input
rlabel metal3 s 99600 85680 99900 85736 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 36288 99600 36344 99900 6 la_oenb[83]
port 483 nsew signal input
rlabel metal3 s 99600 71904 99900 71960 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 86352 100 86408 400 6 la_oenb[85]
port 485 nsew signal input
rlabel metal3 s 100 50736 400 50792 6 la_oenb[86]
port 486 nsew signal input
rlabel metal3 s 99600 24528 99900 24584 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 28224 99600 28280 99900 6 la_oenb[88]
port 488 nsew signal input
rlabel metal3 s 99600 4704 99900 4760 6 la_oenb[89]
port 489 nsew signal input
rlabel metal3 s 100 90384 400 90440 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 14448 100 14504 400 6 la_oenb[90]
port 491 nsew signal input
rlabel metal3 s 100 37968 400 38024 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 63168 100 63224 400 6 la_oenb[92]
port 493 nsew signal input
rlabel metal3 s 99600 85008 99900 85064 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 28224 100 28280 400 6 la_oenb[94]
port 495 nsew signal input
rlabel metal3 s 99600 6048 99900 6104 6 la_oenb[95]
port 496 nsew signal input
rlabel metal3 s 100 98112 400 98168 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 61488 99600 61544 99900 6 la_oenb[97]
port 498 nsew signal input
rlabel metal3 s 100 15120 400 15176 6 la_oenb[98]
port 499 nsew signal input
rlabel metal3 s 100 94752 400 94808 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 4704 99600 4760 99900 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 2224 1538 2384 98422 6 vdd
port 502 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 98422 6 vdd
port 502 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 98422 6 vdd
port 502 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 98422 6 vdd
port 502 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 98422 6 vdd
port 502 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 98422 6 vdd
port 502 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 98422 6 vdd
port 502 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 98422 6 vss
port 503 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 98422 6 vss
port 503 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 98422 6 vss
port 503 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 98422 6 vss
port 503 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 98422 6 vss
port 503 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 98422 6 vss
port 503 nsew ground bidirectional
rlabel metal3 s 99600 30240 99900 30296 6 wb_clk_i
port 504 nsew signal input
rlabel metal3 s 100 89040 400 89096 6 wb_rst_i
port 505 nsew signal input
rlabel metal3 s 100 27552 400 27608 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 42336 99600 42392 99900 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 19152 99600 19208 99900 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal3 s 100 76272 400 76328 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 9744 100 9800 400 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal3 s 100 59136 400 59192 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal3 s 99600 90384 99900 90440 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal3 s 99600 83664 99900 83720 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 69888 100 69944 400 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal3 s 100 6384 400 6440 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal3 s 99600 43680 99900 43736 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal3 s 99600 5376 99900 5432 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 43680 99600 43736 99900 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 74592 99600 74648 99900 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 61824 100 61880 400 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 88368 100 88424 400 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal3 s 99600 33600 99900 33656 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal3 s 100 88368 400 88424 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 59136 100 59192 400 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 11088 100 11144 400 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 12432 99600 12488 99900 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal3 s 99600 70560 99900 70616 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 89040 99600 89096 99900 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 42000 100 42056 400 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 62832 99600 62888 99900 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal3 s 99600 52752 99900 52808 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 83664 100 83720 400 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 60816 99600 60872 99900 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 80304 100 80360 400 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 34272 100 34328 400 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 5040 100 5096 400 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal3 s 99600 6720 99900 6776 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal3 s 99600 35616 99900 35672 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 13776 99600 13832 99900 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal3 s 99600 99792 99900 99848 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal3 s 100 57120 400 57176 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal3 s 100 65184 400 65240 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal3 s 100 9744 400 9800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 4368 100 4424 400 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 22848 100 22904 400 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal3 s 99600 61488 99900 61544 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 60480 100 60536 400 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 55440 99600 55496 99900 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 81312 99600 81368 99900 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal3 s 100 89712 400 89768 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 16464 100 16520 400 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal3 s 99600 68544 99900 68600 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 85008 99600 85064 99900 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal3 s 100 42672 400 42728 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal3 s 99600 87024 99900 87080 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal3 s 99600 38976 99900 39032 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal3 s 100 2352 400 2408 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 73920 99600 73976 99900 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 11760 99600 11816 99900 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 32928 100 32984 400 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal3 s 99600 67200 99900 67256 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 85680 100 85736 400 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal3 s 99600 34944 99900 35000 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal3 s 100 39312 400 39368 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal3 s 99600 8064 99900 8120 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 17136 100 17192 400 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 51408 100 51464 400 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal3 s 99600 48720 99900 48776 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 71904 99600 71960 99900 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal3 s 99600 96432 99900 96488 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal3 s 99600 8736 99900 8792 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 8400 100 8456 400 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal3 s 99600 62160 99900 62216 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 2352 100 2408 400 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal3 s 99600 97776 99900 97832 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 68544 99600 68600 99900 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal3 s 99600 14448 99900 14504 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal3 s 100 11088 400 11144 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal3 s 100 18816 400 18872 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal3 s 100 22176 400 22232 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 69216 100 69272 400 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 0 100 56 400 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 80976 100 81032 400 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal3 s 100 39984 400 40040 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal3 s 100 80304 400 80360 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 22512 99600 22568 99900 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal3 s 100 26208 400 26264 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 21504 100 21560 400 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 7728 100 7784 400 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 48048 99600 48104 99900 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 25200 99600 25256 99900 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 55104 100 55160 400 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 65856 99600 65912 99900 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal3 s 99600 29568 99900 29624 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal3 s 100 61824 400 61880 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal3 s 99600 79296 99900 79352 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 22176 100 22232 400 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 38640 100 38696 400 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal3 s 100 5712 400 5768 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal3 s 99600 75264 99900 75320 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 61152 100 61208 400 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 63840 99600 63896 99900 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 63504 99600 63560 99900 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal3 s 100 90720 400 90776 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 9072 99600 9128 99900 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 72576 100 72632 400 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal3 s 100 20832 400 20888 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal3 s 100 82320 400 82376 6 wbs_stb_i
port 608 nsew signal input
rlabel metal3 s 99600 49392 99900 49448 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3676780
string GDS_FILE /home/proppy/src/github.com/proppy/tiny_user_project/openlane/tiny_user_project/runs/22_11_29_23_55/results/signoff/tiny_user_project.magic.gds
string GDS_START 48106
<< end >>

